PK   6��X��f�>  @�    cirkitFile.json�}�%���4j0�.P���%/��Ҍ1ƶ`<?$� �V���TU[�z�}�}�%���d�I�/�{�n��J��/��`/������w�v�����?���>�������~�����>�����?�����s�9{���>k���k�������-�J5Mfm�g�P��/���٪Vz�v��÷�__�@l�#6.��i6.��6.��Y6.��96.���l\�+��jW�9pԮbs�"x�7�l�`*�+���O�}v_�ܦs�}����7����?_1�H�й�{4�q(.`�20WG����w�����4.�A.�]ﲪ�mV麡���/w��
�G�~� -W��#��+@����t\:� � y���g
0�
0�0�
�G�~� �����
���w�F���/�;b#�*�i�W7Bp�H+��y �!�Dĥ?~?S��� �U	U	�{�Y�%Ϲ#.}�e��V3��^�N���<J竷eV岦TE��Uy��)4q�+n�� �	�]ʽv�����t���j$��B�P�X(onj�sU��#i����>�Q�6�z�?kf��f�;kf��f�;k�.��Sn���WTvu]ՙ�*��PY��6򦨩mu���`z�����S��O1'�hJ��S�\_�����ߣaCx|/��Y�=6�g��maCx�џ�v�?����,��.³���lς��φ�, ��|�i����Y�m'³��N6�gQ2�W�R�h[Ք�QVc3_�x$�gee��.L��~���[�� �!��v�?d�!<�����,�C³�lς;��X+�ܹ�	���76/���YIT��g������w}��Ե�v�gw��qW�gU���&�7
���_���1��:�n �����sN3n�ӓ���
n���݉5����S;K���p��7���!<�/ǆP�\1�8W�ÝΗ�������<���.,³໰��5u��
�+(<8²#,;�#��+;(;²S;�����ʎ����`eg����#,;��X�Y����λNX�9����Ώ�X��X�A����X�X�A���ڕXٕX�A����UX�UX�A��]8�	v�����������/��9�'�N�_ .ttO�8@��#0�p\,?p���G`~�(X~�@ˏ���aQ����
������`��,?�;=�
�_���;|�������=�3�L�\�����GN��L�W\�C������kz��y�R1ŏ�<��<�����/a�����j���؆�������%p�����nX~��b��ݰ��/>�쮎�]O�@�����N��C�7��X͙s�/8p�?�).p����\�>p�STQTu��x.�)���X~�� Z57`�~�|s8`4��:,?�;M�t��p밟G3��8`4��:,?�	��C�(Do)G|�pć�G`~!SX~QH4��%�Ra�Np�STQ8t���>�/Ɵ�Ã���F,?��d���\X~������߈�G`~!�V~4a��_�=�x�ˏ��B֤�骔��ܡۂ���pxу&����/$��/
H.�
�In��̧1E��,xyˏ��BN2���Q����lj`���,?�����G=X~�R����z���/$���ρ�,?�����G=X~����]���/�,��`��_H�x�ˏ��B�?���Y$�i$���`��_Ȁ�8���#0���,?p���G`~!� X~��ˏf��M�%�������K]���/�M����.V5��X짅\�)�����r{љ�T��:4!�b�T�R9=�9:;<���{m�㼝{ߚcI�p�^p�>��e��ʹ9/�T�i�'ف7~� �c�<���t��s�Ŋ.E=��L3o��}- ��܋:&�"n���k���i��͋��/�)��x�А�x��А�x!�А�x)�B,�ۧ7zmt��0m���W}و&:��A2ɐ$F3<K �½�|B0��-��f?����������݌�M���x!Mt���k���_��^�Ԥ՟�@�����ȭ���O�+ղo�z���K�{�Y��/�6���1_�4��zC���ap��=_3/��K�Y}�_Rn1�P�I�i�4�5�:Y�y���U��g�=�5����\�K�A�0]����]�:
l������ܹL)�ꢮ��)�FIՙo_���^�e'����H����$U_vv��/;�I՗�4��Sx�Լ3�vZ�e�K̗ċ����T�~�^���9���(R"���@��rg<շވ�*3Uc�r�6�3�8��r�h�Z�T���]�٪k���L���T��ƞy{R���4�W��TSfK����͠�2ﻡ"��3oO�~���%mfM��rUV}￥���֮2չ��T?#���\[uYcO~(}�����U�j�W��=����_����������>���R���?���1$�
�aR�p`��Tp�0�@@*�WF  \6#�
^ �H������aR���0�ѣ�H��ƙ������29���/]��LN �q�#C�[�<���I��톡e]N0�q��#�چ+'�8u7~]��I�!�~W��̈� �`f����av���4Z�JM���@Hj\��I���d}�&'�8=��/�I��-���~�k@<s�H}��qҸP��q�7�av\��Q(�i`�����換���-J��@H�6�QN�;�LN ����v����(���	6�b`v����8�츁�qR�
�Ą�q��(�pX�	6#naS�(�p�	f�-̎��B�>'��0;�B�n���PH!GLN0;�`v�r��8�츃�qR�y����0Ҕ%�i����=�Bw�������r!���0�5 R���q�?�`v�4��Hu�
�]0!��*�E|��av|	i�f�i�8�	�J"\I���M���Q�r��J"\�n���
��W�vӔ�pT�\%��Ww��u��#	�$���A"r�&*�H@�+�p�>��\�	L1��J"\�n���
��W�v�T�pT�\%��W���@���*��D��=�2��L�%d؆��2��#�x��B
�d�.�	�H&�aK2l�^s��D_"lI�m�3/#[�L�-ɰ{�ed+���%����le"1�$�6�Ő�m�@��pl�-D2�QD�2!�[�d�2�#�le²�!h��LǑB�"li�-D2q��YaK2lÙ+�ƑDo���d�2-�i��L�-ɰg�dd+���%��,_�6>�ǃE�V&.a�$��m�@�L\6�"��l�%[��l�-Dq��	2+e3lѰH���eZ&.aKslB02q��Y/aK2l��c�ʬ����9�!��eFf�L�-ɰg�ed+�[Qh��L\fd�2#���%��W�!eG:{+�Ͱ�!�t���Y/�a��E�V&.32�Eؒې�AF�2q�[�arW��Vf�[�arp�����e"lI�m�%"#[��2�$�6���'X��l�-)[�����e"lI���u�H�Ƒ"vaKsl!B��ˬ�z�[�ar��V&.aK2lC�#���e"lI�m��$#[��L�-ɰ��dd+���%�!���l�L\&d؆�`2����Dؒې�LF�2q�[�ar���V&.aK2lC�9�ʬ���%�!w��l��|����˜L\�d�2�$�6�2���L\&d؆��2����Dؒې[RF�2q�[�c˟92Ed���e"lI�m��)#[��l�-�d؆��"�e���2�����������v:+����C��E�g���ܸ��Mw��9�0�e�M�ވ2f���8oD9���.oDY�Aa#���ј�:�F���W�WEeW�U��*��PY��6򦨩mu隃��Q�ڈ��}x#�S���=LQF}�o�zE��jJ�(��������v�gee��.L��~]�I(��7�,�}�ŬY�$�f�PܚeHB{c|�F��[>^Q
�M��!T�2��.���f���*}���nᾉ�(�������P�ZHB��U띄�p��F��,��߈����ց����pE�V���$f��H�Y�si+��5I[a0:|���ܐ�S��iVO�Mi0�懧��5W1f���&׭0���n��h�^�D}+L�6���<��ahsLuh���6K�n�Y��}W��B=[�H��uV��eJiWu]TM���$�`��z5I(��:($����$��!!	euDHBY�j�PV��4�)/F{	�����u�&fU�m�UNg�.��-��(�5�*
]���˄X;�0nG7�oDY���B�:˝�(�o��UUf��{�C_�9���$�U�k�Z�T���]��ۮ�ʺ+2E�jSi���%	e��1MC}5��5e�T:�:/]U�y��\�sIBY�b�PR�fք�*We������m�|���%e��ʪrm�e���o�Y[١�[��*A_�P���2������������+���������}}{�o�=e  5~+�H����F_��F�	��F��F��F���F?��F����/�D�6�l��6�7
I�|'��&��F!�C ����3�($u���p��p�q�:LEc8�츆�q�:L�c8��o���f�QH�����f�QH�J����f�QH�~����f�QH갲�	�av���8
)d��q�ͤ�R`v���8
)d�q��q��(����	f�̎��Bf5'��0;�B
��`�`v���8
)d��q�͉�&�av���8
)d��q��q��(��Q�	f�-̎��B��̎;�G!��0N0;�`v�24�8�V7q˛0;�`v�N��8�츃�qR8����9̎���Ia'��av|	i����T9�p8�J"\I���E'�Ѩ@�Jp%�j�&G��*��D��]���
��W���.�Fɽ ��J"\�$"�(�D\I���QD�%��H@�+�pU�(�(W	�$�U�l^hT�\%��W��2y�Q�r��J"\Þ`��@&�aK2l��f�
E]Ba�L�E2��D^"lI�m�k.#[��K�-ɰ{�ed+���%�aￌle�0�$�6�a���L$&d؆�2����Dؒ�p�DF�2�[�a����V&*aK2l�����L�-ɰg�dd+���%��̕�l�VĄ��d�2-�i��L�-ɰg�dd+���%��,��le�2�$�6�I���L\&d؆��2����Dؒ�pFTF�2q�[�aκ��V&.aK2lÙ]��I2q�[�a���V&.aK2l�j���e"lI�m8.#[�݊B�e�2#���L�-ɰg�ed+���%�!ǀ�le�2�$�6�J���L\&d؆�2����Dؒې�BF�2q�[�arp�����e"lI�m�%"#[��L�-ɰ9Qdd+���%�!���le�2�$�6䨑���I2��d2q���ˬL\&d؆�A2����Dؒې�HF�2q�[�ar8��V&.aK2lC.*���e"lI�mȩ%"['���%�!7��le�2�$�6�8���L\&d؆\m2����DؒېsNF�2q�[�ar���V(ˇP������eN&.aK2lC.C���e"lI�m��(#[��L�-ɰ�%ed+���%�!G��ls��L�-ɰ�>ed+���%�!g��le�2�����������v:+����C��E�g���ܸ��M�t�F��ܴQ��nDY��e!��F��\�Q�[oDY�G�����꺪=@SeV*�\�fC�5��.]��/I(������/I(������/�UM�e�16�]�����L�ׅ)\ݯK7	eU�I(��MBY�n
F���1	e�7&����BkӸ|�U��v�˪��Y��ʪϛ�\ח$�U}IBY՗$�U}IBY՗$�U}IBY՗$��,��߈����ց���KWvo�������[a0�t��V�/]���KW)o��`�/�1���K7�n��h��}�[a0Z�t+��Q��Kw����]�:
�l�#]��Y�;�)�]]�uQ5źW����ڡ�PV�S�jwJBY�MI(��)	e�/%��v�$�՞��u ��h�W����u�&f=�봡��l �eֶeV岦TE��UyB씄�k���6��T�_g�3E������L�آ���i���PV��jUS���v��o�&+��Y�M��o�:�$�U.�4����֔�R��tUY�}7T�s��%	e��5CIE�Y��\��C���+7�������6*�ʵU�5f�_4���[fme�*o��}IB9��˵��_}����~w����]_�ts�?�>��m��n�v����������y�]G�Z�]�<���ڬ��_���*��2�}��sƛ�w�y�c���^�WΫ+֫5G���j�|u�z��|5-�:q>��Ջ�+q����Ε�"q���͜���7��غ� ��)Z�}�5ʏ��3��V�DC����� �����e��'.�\��9�͆�നn��8��/v�����y�g�W׉eX��|����0��~S��#���\��Ԗ�C��L�-�:�˷7L����Ǽ��*�A%�3Cw�q�8����C�p�Ļ�8Tr�3R�>g�߯	�ĸ��w^X���xg4l^c� oVE3߾�n*.x��;�}�シ/��
�`)$I>@�f�2*���z��rl�n�X���"֎���Bt��o���� )u/��!J����V2R�0��f~
3ؔ?}l�f�9�L�X��@Ml�%1E��>Jd�29���er
"�G�����斃z"�[6s��9[�� �-noO�[d�!������/���D�w�s_���z�)͚��/���a�0N/Xc6�f��1��L����3H��Q3g���f�$�c����ά�2`���5�C���0������t���6q���L��5U�y�6��6��6�&��DXρ9�3�W�K�oM�'�6V�l�s�a�<:%�k�4LiS�i'FxzS
:����p����ڄ�o?�
u�����=���rvWh�����~��l?��ɘC���\�w��۱�_�Ts���5o��G��?��������v�]7w��[O����>��E�{��π{��π{��π{̊π�u�π{��,�79{�g�=��g�<��'��N<�|o��,����px��a�Rw��m��8-�' 84�'8;�'8B�'�=I��e�F�m|�Y+��'ۘb`��(10�؉���DF��#�$6��F��X���4��6�������ϔ�f��yG/I̱�sL>H�������'�x�0O ���-�u���ޢ�A�oQ!u���7��?G�M���7��cK�;� {�̀=����6�����?$�Wb�ث�l�Ğ�c��st�������|�:��:��:��:�?�Fg��3$��@��3��� d���\� �O��������d��$���ȁA��d́�`'�������������f�9k�?KR>#tn>#@��=Cdځ�-;��M yw�$ �w�$ Yx�,I���8���.���3+L\|I03�$��q��~��I|F�I|F��I|�,J�E$S��T����J�K�F�'Z°B�[��"�� �� 	� � %�"3� A� O� ]� k� y� �� �� �7�� ŀ�SI;>�8<#@<�A%t�.@�C�5���"�e��9�0�Щ�0����O���j���/Z��YҬ	��[ת`A77�@����j՛�`_�~,��&d��;y�`���g3��N7荀�s ��s�ƕ����n�{x���/?������~�馻��3�}�C�x�$>6�� >6�� >6��Y>6��9>6���|l�+�,�jW�Y�!Ԯ�`Cx�0�|�qr��#`��?��r�1$V9z�$w�9z�$s�94SH��r����;��������iqcV� 0bLh1|`D1&��b4`�1&��A���={Kr\4�/0xkQ�$\�����gP#H�*2�4���Z0
�� ��!��j&�� 1����� 
4`�3c S�̌����4����9���`s�+�!ǽ�$sm�Y&q�a�=�`� �:�� �q>�������p�1���u>��0�|�p �0#nS�|�p�`O-���1<�=�c�p8��`Om�s�����%���1���-�� X[>����|�`m�c��H��{��c
�)�bnW�C�)B"H�7rL!A2�*8�g	������1Ƅ@����z���%���1B�D �c�,u�m��s1�̏��Ԏ��#�����O�4X~,?,?�S;���ˏ��|���ˏ�������ˏ��� �_�����]�_�����]	�_	�����]�_�������h�����A~�#/�47�l�`�4C�+t\B��̐�Îj���	�!����h�0CB3���2D)`��f�ʣe�T�	��4iF�Q0p:Lk�0`�4C�+t�2M�q�|�@�31a���4����H �Ą�s��g�[����&��!OL�+tȣ�/`��fx��#�(���%+��	�a��!�F�<`��fN,�e�y�	�0�;}�`#Rtfx�`��Q|1i#V�:B��\	��i��hޒ�j�	�a���b"�]���bD������4�@�(&��d��z�̐�O3�ad���Ü� ��\	�"�^�3$4�p"-C��4��4td��AG@`��fxz�F�Q@1qי�%�0��J 
(&`���$bD���z��!����h�c0CB3'��2D�c3$4Ð5 ,C�j�	�0d<@���fHh�����0�L�m�AML�):���̐�O���0
&z�\m��\	�c�^�3$4Ð�-CtfHh�!�
Z��(̐�C���Q�!���6h��0CB3�x�2t�(̐�C&!��Q�!��,Hh��0CB3��2D�-`��f�O�e�^�3$4Ð-Cx� x� t���q�C�)`��f�e��S�	�0d=C����a�؆�!:N3����u���($��4G�-`��fR�e�[b�-b�{Y�V3o��WN�(�Z��gα��_�J��y9���J�"��Pee��Y��27��k���䑧I^7��w\�fc�_Fq�6u#���
\��|c��Ե�t'���u��d�7g+*���j��T�Յ�*��ِ7EMm�K��).V4Z��$�(I����fтf%�ͤ^^�۪�t����y�a�5qyVV�������d�p-}\��uc��+f4n�W/؜$�X�K6'	n��/hF��EY�?	.J���(����gT)�qf��YP�$��YM��ftg��&�����՝(����Q:�V^����лd���҇�4�3N@tq�V��Ɠ� \-��uixIË/�[�,�L����*oƳ�ذ�KE���4�X�5�(�]�ɱ��-�[֮Gފ;�K.C^�!KA�a8�����Y�Zuj�҇�.��2w.zꢮ��)�9EI���?�%�7��gF���gzPR�3cFR�3CFR�3�MR�3�M�������UA���9�%���N���R]fm[f�Q.kJU�p]��3A�Y��H���2|��&�ţ�Y��P���x8շ�\�*3Uc�r�6�s&/���k�Z�T���]��خ�ʺ+2E�jSi�{��I�ϼߘ���|��2[*�U��*˼t�Ͻ?����[3�T��5��UY=�����rC[;ϟ}J�s�/�ʵU�5f���ҷ_aˬ��P��}u���������k��n���y���?_�LY^}��*��=�(>x9���aUq���U���<���2���"�Y��
�a�FF}����Fo�_gEǠr��|9cb��z���ql�yǔxc��1��s�=�l���#O?ł���'X����J)v絒��b(N*����
	]�սnm�f����ֽ�d�&\Y�-ˡ�ޗt��{K�s1^���7��oi��[�{���)��]�=qw���t*T�|����#;֙�x�1f�9�Y��eg8��P�eg�%.qAW�cv��E�^_^�&�7�'�f}bi䜶bf���̶r��7Y���eq��V,ɒ+ɜ)I��r�g��H��J�y�����g�g}�Ē$ŕ�eJr!�OܤÚϏ���%�&`�Cӓ�1�%(qs��]'�05����Z�]Լ������/�2��X���$�te�:)f�8�)(���bv9S���i�Y.�H���cip�����.�Ƃ�����k �χy�y�;ͣ3��F!�5��[����sh�ϡy�����]��0�zy��<#�3p�u��0�>�$bԌD��1�?�*o��/2�nL�n��O:u�F�E�~L�~��R�|��~ӕ��(�8�;y#���ϸ����a��k��r2}��L1C�/�׌Lo���|��.و�|�pg�a���,ř�[Ax:X�x�f)�L�
�c�&;��Թ����!��O-���c����m���a�UM�\}��]��.(��	==���~z��G�鑉٧G6~���Q��(�O���Q����UO���=K�bqЋ8byг<(=�b�гD(	=��b�гL(
=�b�гT(=��b��g��X.�Y.:��~�v�~�c.��}&~�y~���g�����`^s�ˋ>���s鸍�s鸍�s鸍�s鸍���L�>��>3����q��g.��.Է��#us7�w�7�����)Ⱥ:k��;�E�d���?�j�U-�;��u}����B�2�n��c؝�b�r�k������6_�Z*{��ĉ��2�=�s�X{���_}s����?����?ޅ���E��xs�g�=w��������/���Wb>��xrW�_?����������>���y�in����������><z��~��>u��龿?���b�,~�������w���>�:�C��<-��<��<�-K�^��.���{��y��
�k�M�x��\��P�/���}F��3=�0lp�u�P���]5ȟ����Et}us��Xߵ��Mr�W{��w����U��)�R{s���OM�mQ���'�5U��������b��i��RF�?�����ص���S�<��x}�?�r�G�ѣ�V���<�]�<���	����Q�y����O���E�W�޼7��t�I�Wth�g�rm��\U���6/�7	eWd���L�v�T�ʬ뚎ڶ�f��ms=i���6����6�6�z�PuhLWE�d�A�T=���=V*��K��xj��Gn,^T����x�
��<'/N@s�Que����{��֖O�s�Z֫�s&�+�M6�L���:3X�S�u��zh��ik�������"z�/��IT�T^U׾K�/��E�V�:��JZxy�*��o�Jim�ϥ�U���V!���{����ƽ�2���6�,��o��&3E������}��ρ*�7�V�C��L����x17t����
Cemᆬ'���-E6�/�ks=:��*��97Me�-�DcUУ�#sY���C�ps�|�`��S�K�zi.�^�����IK�F�6�X��C}���\]{�W���;7���� ��������'�4�>�y-��=��(?)>�[��h~�����O�u�������(Y�ۿ��c�߿������{8�oZ���	I{����*���u6q*����j���;0a˔�o�k���ݢ-[W'�p�~�����[�t���N����ʹb)��菞�S�\⨅�tb"=x��8}����o�p���Vm�Y�ۛ�_?7�77��<���˻�J�MS��������������辒��y���?�?����?���Ͻ���k�,|�+Z��������g=���x���,���W�jm����O�#ܿ�]��9z������]NT�.̵w��;gs�))�7��ɺR��Ym�*��K_�,���m�ՐԷ�Nj���7������M;g��/�Jʩ���M?d[��0C��RWƉtͤ�QB]sK��1Nɿ���W�ݧ��=<x��ɼ��}�p�T�*�M�8�LV��e�7�J{����{�?I��[�E�o�ֶ|_��/�r���X�U-�2j���˵�r-�\�\~T����,��Gz��]���Z�F�/�5�t�V��#s�L��g�L=w�^^-R)�YV��-�2z������(_��qۨ՗��h�L�9m�+6�s�f�d�X�1��A7�!N_�ۮ�������}w�ừ�������������-F����:+)L]��1ރl����������_��͡�-�̫�͊�k|�VgM_h�*?�)ݏu���꙼1M5tYQ�uf����S�3C����{�������*;���Z��ʛ3�^ZdU�R�M���P���7w��o�L�{�ׯ_��7��1-G]����&�¨�jl����v5�y"��������?�w���Ն�2L0�̚�����̨�X��nK4������?f㺚
��0|�1��:�"+�nh���s�?}���c}�����`~wU�����ԯ����~������Ow���q��=k��o�����������/���]7���r��y�~R0�jԹ'�&�y�E�.�h��O�˺ZR0�?�U�٦s��eu�t��V5����fN�]tu5Pֵ^3lkˬ�;����ڦ�+��
�ʰhS����iq]k�8/x���ޙ�<�`���������=�>������ﾻ{����ݻ�yo���](�����~��w������|i��/���@���<Ώ����}������o�`��o��qT��x�{���oa��7S��dZ��}����C/�L�����2LJ֐0eh�q�p���>�Zx�騕��k�!�=�$:����SG?�4�9m>m�{?ʒy^�(���I����;�9Y/U�63>���NSg΄�NW+�{��(�5��$���c�yīn��U�������EsW��e�0S����_U=�;{jP<ꥒ�����c�>pQ�ZU>��}λ�UQ����N�H��>o͐5λL^ɼ�x]�F��s�uF�;���.)]O��wb��ٰ:��o�/h�'<�:}V���}P��J��4g
���ѫ�8~R=��-�i}\�AL�B�� �}��r���ʱ�jaJ��������0��N�{�}n̂��ǁ7�7�Ge/=�^�C+}�FCS�>$4Y��vN�G�����m�h(�$5JJ��e�������M�Ǭ�5���a1�Э�^�W>�w���7�B�wO;���~����0��������[��t�m��T��)|�7X�?��W/{W�����������m9ڳ�C��1���_�:|�8z)�?~ss�*_�����u3P�dh#�}���\=޿�����{��~�a��wWa3��o?�=�!��÷��Ô������C���Ix�Xʝ8�/��h�\������o������,Ru��������T�g�L�	�)sJq<L&�r�fU���T���m�*X�l�`�`�ty
6.�ͨN~����>6B/�rsj��J}6��)ނ�
�`f~X�'͝Vʙ��/���$,XZ�O��хlW����ݨ`��fvG'���p���&�).5�:u�r^u.I�zF}��S]ӖWz�ç&��p��g~׍��ʓ>o�Y�0U��R'gq^K�+��LU�yU�X��E%�K�%�c��8���)��4��|ɢ��R���[X�4�N�!�R㶩؟9�:S
��宆� �T�`���e� ��5����}�S�5.5�:��a��>�;��nM�-烸���g�w���^��3>HT��TE�W��5OdTZW�*B|�y��� Q�/��7�! ��X�,��o`��x�-�Ը|��K}yIڽ���T�E\�$E�-8-�� ��d �Xʜ�*WJ�+�З����%m�<� (�{&�?Sτ��=�J��AY�L�Ro�*꼪\�y2cժ��T�̫��3�J})��N��ώ\��:������xm�3�J}yI�=J���z&���ĥ$�R/Y�NKM}�m���R�J�y�j�6�B��r�z��B9�gB ��T)�ij���mK��z3UQ�U�b͓�VՅ���dA-&�I\�Ki��w܉�6xΤx&l�t{eR��l��g�����{	E�z&�M��$[pZ�%��i��ϱ���9��ԂB5e�wu�m��z/��BY�gr��2�L�y�t2E�ެy���X[dƗ�&f�ě�o�7��6��ZE[<�qQ�1�&��PJ�����{Q)�NԴ{s��@�kt�w�l�
<�1G��D'�͉K6��]D�mn{ᦟ\��=C���'���m�&�sz�&.5�:���!��hK\�!��خ	��+�M�U���z��U��bmq֛��>7q��'n����/Bmm��X �ą6zrn.��=9^��&N��J�	�7G��P�;�M���$8�M���2k�f�ؗ��_��!�7��,5�d�_j�y;2Y�O+��6�ܔ����/p7pF<sty-���WJ�$��݅���枡{As���䎬��5�PJN��آ��'8�5��F6���v�Ӄ�\y��K١�\�労�(��*��Л��:�&k��+��*,5D���:1q\�B_Jso�� ���}���ͫ��Bfv����)������:�Y�Z8�l��{0�s�6�w��ƀ�"���<eKFZ��;=O��׻?�Bo�&꼚\�u2�iUUXj���ub2E�����j�e�<]d&C�|��!#����ɦg�S
���W��(*uq0��(hd.���~S@}�QЫ'h0�V�)Y�����x������n�CV�q1�
0��c2��Z�K���w�k��A-�yPnԘ̓YR
��ԗ��G;'��;��^$e�G:W�:�Bj���O܆R�7������`c-�oj��Bcb�l>���'&�|�ߺ�)����YDt����\Pj�Ts}E5*��ʂ�8$�,��CeYXC5��*K���BO��sk�%�>	%�Jh>;�t,��})M���I����F�a���y��b�E��"*���b�Ik�����"�EϏ�Z�T�*J�s�M�D�)�H0eaR6�{���]�o��[;�l{���E�N��da����)�,DTjI]����ꂝ�$���+	4_��G�hoyT�Ki�N����;#��,5��XIj1��rK)�&.�4��~�;O*�.O���'��[�"k�R�|kLoM�RDz�&֧��R�!��N9���W��t}�άN��ǒRIp�1a6?]��nm7 �l�!��7ڀC�Sk���z~��tN\�-�`a�v�m�Q2f�W��c�3U�r�k��R���z+X�1Ő�@Rbo9T؁`ۅ]�����wE*0��1R���[���e��X��
�.�c�sU`>�x�Q��T���^��[���]K�\��'R��"__�&E�P^��/�+r䟡���u��K٦-�� I�� a�Q��+R+�f@��RT�"wV+&��ߊb��:b�F�VN�p��󆋔����o��P�j��L͑�5�������)���jnno?��~��o�ۇ�A#�n���~[�}�o�������Ǉ@���5����o��h�o>>���|ū_�/PK   6��XG�~��  � /   images/0739a1b1-a163-452a-a325-ab452d55b136.png�y8�m?�r�J�M!*IY��Ie�^Y&������[�d�cb�0��d�1̒,�ٲ�L������������|�|�4}��>�r}��|��mn$�_l��mۄ�o^�ܶM�i۶]&{w-�����A���{����� ��n�m�&�I����em4�6�l����
�*y�����x(����WŶm;����5��9t4Gb&��Ȳѹ�}��OܜΉSٱ������b��MT�}�L�1HƸD���?j��i͘�ǰf�	�A��{�ξ�[_����J�z���r���٢w��/5a��t�I��ե�EnhǶ-?����'m�ں-��Ǔ[�n�-��v<����xN��J�h���e3��2������7��=V��)u!";G?�� ��<�|K0�yY���I2,���^)�Ϭ���Ev�p�����������d���4���dK;!-�L�^�$Cx�䐦W��k��E���9謗	* P��ϕ�����S�����0C���~�?��$Ǖ���φ%mXJ����{���w/�y|
�T!��;��G����쳄�[�����⩧�U�6}3���6��{�[$��ab1�P��~z�3������Y�q(�V�f��¦�&	�� ��l.Z��s9�2SH�W�ơP6�[��SnT�QokF!s�Ǔ`��� 6rl�������fI�:�v�K�|l��%����)�m����}gw0�6=y�dk��?�/������<�w�}l��جJ���s�+����������6����Í�͍{3�����"R-33�	a\yoU+����̡-�߶~�S���v�ѯ�f��nY7�߼�K�pE߬�����f�J�\t���+"D�,�����AGf�H��X��i���&���oց���A{10�^���l����UL&0���ٵ?���E�)�Q�5��s�=[�,�8�v�Y����>\��>\+sS�N��88y��</�!-Ot�HS�/'9��q�ZwuR��
���ӝ�v�����xS>edf5�Ի`��Z��/�j�3�QM�/
�1Q �wH����G�h�p���"[�|���fi�h.��-
��f�:�[<?>gh8)�2d����q���j�GZl��Ϩ�4.{��F���Hq���5�1͸�m2�2~�l����]I���J�&k�-�x�T�/�O�z�5�k����8��JdX��a9�<��V��\�����R��9�����0�TƦ%r�hm�[o���b�Pԓ��YپQ5Y�� �>[Զ�f�UG~����bhA�A	���6��,-��:[��Y����p���m���k���A��p�ʂ�K��&�{sdJ;?=3�O�	}�Ij�>>wE�Ws20NJ]=X�uq�g�j����bN���|�G����Q�s˪�r���W��ӕ������7�[����v�ЂF�K^��FY�{��s��ʻ��R�:i��D{��x�����T�Dr��j�M�s3�����:u˙��[�.�[Im}�v8��0��d�Y�S�ܷ�BW�V�F��V�E��V�
���355;����҈�RW&/�+�'��]W�e����v�@$�Y��=�Vܲܽ��ٳ�6�tinb��[s!ޞ�C����<_��iG�Gn���_a+*�� ]>��-u��{\lrǹ��x�|�b�ߕ��?e��@�㕸�����[�`J�p-��i��m�'���n��:l�xm�pd�l�em,W0Q�:��"�A�fXDyP��pOTG^uPiN��c��+l����~ŭdyώ�ȂrZ�����?���A�Xc|O���/�Pc���>���tx/��g�N8^xai=���
\�ΟNXi��@�l��]Q�0��!a�+ץ���q�����`Vq,�o"�B8a�i���Itq�����1C�06�J��J���
�<-VTy�����kQ
�ɍ������p�F����Ϝ����r�}��O��u�~�Ar�u�����Wc~2�ƪ����@�m�����
&�H�;7��.2g�>)l!�(�|�v�z��[�TJ�й��#�J�:F���R���:oȼ�>33�w��vå"����P|�?{�&��#�H��+���#��<o��Jڐ(-�������&�Mt^��R��|٢����q`�g��c��j��02���)����F�;W������+�xR��:P��/�ސc�H���\k�Ý�/���d�����^� u �Ƚ���c��������-6yK�.�d�j��܉�x�������7�.{��"�'�>����K�۰o�g����m%���UY�> �/��
zo��X{_�v��Kû��q��Ŧ�ү2#G�_Z&�k3��x��r��2#zל���@�[��װ��^_�L�#/=lql�X4Xm������nq�p�7ME]�A��J60��e��ogU.Ė�FՄ�W_Ћ�[cT���l�hze< &��x����/{�"�Lv��
��= з$:��Ln�_�|_�!��ɬK{U���G��Jak�6����������R3Ć��S�ۿE$��|��ӝ1��E}��q[s<w�R��.�$����V�P���Lկ�0e�YK�9��qO_L���p��Tu��/8�ˊ��Z��]��A�@(�^�1���s�z��'�l��x�}u��A���<�� m������j��1õ��B��iB��	�A&q��6�t���+�cQ"M	��յN�I/&�'9�˹��Vv�t�R��FAD�/��"������N��+�',��Z.����xT�;(a��C��?����Drɴ��J@a��m�e��h?-����b	���M8=�^����=�ӽ�b/��Y:#�3���rp`��$G7��0_��s�N���vo���B��
]\�R�	�e�1cٝ)z)A���۹����E;DO�V$���t+˾C��@;�sA����.���8yQ\��Gwz�O/9s>u��ř����e�5o��e=���qפkx�t������]�o�O��V��f(�\z/�x�@P�p8��R��fU�j�nL�`v\�\fM����qY�cGr�?�������@�W����:��7[�zȏ����{�N�ND�v�bKT�
{���=��s,�{B-#+�Vx�Z�%��/�(?��9&s4]���5���3\>�P(y
�6*���+����&�sN}wT�$�8���/Aa�ԥ5i[����x@�� �`��������4�nc��,��R���1��q��a��­��[C���	�~n���7a�F��G�S̻1[�#ݹ rŀ�}�uNʂj*�6I�VU˕��UP�����h�1G�2�Rs���Ծ�y[�J�梵3d������A���i(Β�����~\@?�,�8�(ݙ"�i��ݤ�܇^��g�ms*$��ESפ�#-
!���U	�����lQ�̵��K�1u)�ױ~Q ���16������	���8@qY�&C��.:!�6��;c0߷s� ��g��"HSK�P
��10ڂ�|���}��([��`�d>�*��I6�c)<���H[Y�ғ���,~ �lvЧ%	Y�m�[��>+�8U�t�@�e@��v�AB�a������m����p��_ \�**�>j۪��q�E'|���s��}��)��Һ���w,���n�b*� M���1?VPg�>V{���M�|j�:`�@�������x��Ox6���Q���s5��I�a��P��'��C��ݽ��(��/(���Y�<x�̶H|�d��kѺ>�Y�G`���*"�r��l��$-.���A@<��E��u�#�n�����,�=�bB�B��^ͧځ[�<C��^� ��|�C$S+��G���.Ԟ�*��� AP�	�oe���W�\t ��i����� �D=CZ7��<���?��1����m!�����;ZЮ��|�-����;����ٱ��rO"���_�yF�
�`��!�;��U��X���t��(�JW9�~�#&�M���j�n �I=�x)��s�Y��rvHYF|>zBf�؉P�":�m��'(����n�?0 �捻Dr��Ox@{٭�Qh�BU��_FQ��(p��
�zk6=U�E��+��2p����v�)��Y��4`�n}��Ƕ��.E�Tes��q�e� p3I�k	Y�պ��ľ̫�}�Q�@�i���u��<��mЭ�6�e@x~_�"^X��$Ԥ����txY��&��_�/薳�q�1:z�3#9�Sd��V������#�����m8./����V+}����� ��jm�*~Ԉ`*P�,��\aK ������=}�������1�c,��s��E��J��3�2doR0�e��&��}
�)@h��}�G,;�`�͉BJ�Q��ib�]M%�%ᖝ�$�3���0f����9��.����l�O�u+6��,w\μ���� j";+k�Q@��7�HDi;w��d�N�Ž�͊�BX���+z���I��Ӎ�R��2��q�:�r��Ť ꛕ�4�J�\Dt��>w&�����Q�)�,m�k�b��	�KM�PA9A����C�T}�v�٥M���dҊ-"�Ҧ�^���o"�.��Jf���Q�^#��B6��&���(t�f�4��g~yŪ�Y5����A�Epq�3���Ĕ'�Д��*�AT:Vb��|���-%�uw�e�I��UU<��2Pl�SF�׋���t���ޝCɶ]+�7���Ld=>e�_�T{�+�F^Tx'M����DE�o�-l���P�G>���Ѐ]
�?�8a\I��$��B�Aِ�"�n��P�j�����Oy��eDH��t�k#�AX_�&��O�-���T`g��JK�7J��"�Ÿ�(64U��]'�YP��D���я���rZ~�xy���uu$|�2���d~���a�sa�w/���������&���5#k��'+��}PkH,h�d��v���Tϴz��Z��G�_ZN�ad$	c���Tx�4�nʤ��6�P�����ʞ���|�uxP�[�+l��VF�߃)��k�~1s��Q��"���c&�,�Ƶ�ͦ�X���ϠoC��l�I�v�$Fc�I��2!cY����RI����-䋴X�Za+K�k��Z��\�=�Y����n4a��gT���SQM����܁G�"�]������ ��wl�q-��/\y�u��f�ň7'�
�l6:�9��#�!X�Ě��b�����F����w�:N[h�[�n���=��C1;����M9"〧����;/Quu������� ��N�ۖ^$b����|7���V�Â��a��s�.X[�H��M�K/�evTv>�U۟��gSǄ�E�|���Hr2���}U{9��y,{�hh����y� h9��&5�Pg��X�s2� �b��ͼ�tzer��;�4O�+NfpE/�ݔ��(BW��r���9����(�oB6������픴Lq�K���xRtJ�?K((2�~^>��npM��Y��#�)a��ݡ"�#�|�a�*�*�j���[e�G(>�D/��(�|y�W^ x�m#�]���h��0T[fLL�j�~Ԅ�jo�u��9���p���r~��So��}�'�ť5^LP�1��
IJ�p�C2�����IJWC&� ���/��\���=%ݰ�){�����{8�ގIR�v
�Hp*Mi֪�X;����SAe���x$��V+<�$���s��\~�z�}x_a{�x{���#2'ͳRl"�/=?�z`��V��s����8�>�ȷ��k��*98��е��zy�i��S�h�4�?_�\;���Yմ%�V%��b?�����ܕɪq�ꑝLO�t���RT�^d.��p�*�> '����'b�CU/$mް�Q�ql�[�3@��pu��ToV�@���Wz$�jIgg.��]bT��$%
�?�H��4(eh��Խd�,�m��cn��B��
�b�9�uLT3��	yX��a�*O��;۬&����Ⱥ�6Kо�S��`�\�˙o�
��Z�d���%�����隲��/�@,���z��҈��I��cW��f�HЈc���h�|���Z#��Rt�Kj��N�\%�����n{(�ډ<��3�r��AI��֞��C����Gz�.Zm���J\i/��I��)�k|�c����l3	]݄K����'�q#��+��?_v}c�1N(��ߡ��~5�(5�T�Ӥ�O�!��n���0{HMWǥ<�����e��ؘ298���i���|IT�VDb�*y�>w����$�Om�~W�z�n�W(���r�
�z��Kȯ���'�q?Z�X���U/7���3c�n���e�����հ���e��Ym����� DQ� &5��}z)t�ȩԻK����k<�q<�2�1���<79��������8��в��u�F�'Z{r��(ഏ�,5O�o�ܙ�v�ʨ���Sn)ړ	h:ͽRj����D��j<s���Y�H�5R��z=�B���㼌��a�}���UZ�6�@d5�b��	��sV��5�n��7n�:�m��!�'u�	l��1*�Pte�
(���l��U��<$u�{�<l��F@�O���Wyl�@�+,�)����a�
e��k���O�X3��J{n6�Z���G�6o\�]ʚ>��R�,�g.����{Y��ma
/0���U�υWcnI�*%\��W�+�V�`õ�x�����b"�r�=�\����Kmk�)3��g3���	Y{�D�}<�76+7Ŭ柕� o�|feQFW�C�:?��\lS������[7tُ`@?����چ���� }zY��E=	)?YQQ��-ח�q��syBk�S�3Q�0�w����`�ӷ��FI�e�c�B�g�Y���_���x��l� ������l�MҦd� v��q�P�>@_�����^ZiE>�)>���K=��*�ڍI�t/��.%S�B@�����T ��/��GJ�{�fm^ͥy8��ro�Vö�ϿNo����i���ѓ׹F4�6�>jY�::�zֈ�K8�Ϩ]U5�SX��k�<����)�Q_���ߙ�%���sY���}�Q��*��4f�d�Q��*VE�z�5�
xI##:@�t�}��+�{�;��$Mr�J�������/�\��1x��U1y(¦}]ĤwD~���C���ڣ�1��H{�g�d��4=�Qa���M��QZ���ը��fGR�}�\��8Ғ�q��}�4;l��/LoF#�T��7����֍1�ޣ���'-�xT�C��h*��-'�I��M�ڈ�s��/�_�{�����G��L��z�����,�+����F*�޳V�����>S���D�Rg����;�m�.V<�����3�t�`#����N������M1��nܩ�7��u&�]�{جʦXO�k�௛:Rg�L2�4�Z��O�TS���q֟[� ���]�h���uj����X|��Vmwa�O��D�����K6}���n�Z��Oe��b�u��2��A�:vq��L�J�� C"<��Z��������������;��X���H���[���jB?�ݧ�#��Lr
���-T:�+�D֗��@�E�ѣģ�|Qgp=��F�uK�ܫN���Q��� B���Ƽe{\[7ҵ��H���n5֎6�~�b�.bצ�!�P�	�	G���k�눸������J�|������^B�^�Y�n����5��f]$g�(M,���D�h�t`&ȍ�f�j�7���xYg]�22X_7�����=��f��7*qKn�ֱhUr�Y�}$U��G�e��_~�T�1�;��j&�>��!��I�.�*۬�=��(��0T�	�GU�Weh�7bTQ=5�8�n��މh�\�_����+D��YZ�wr��V1Mw^im�G��@S�ɚ��� �w\E���Y�wStH���n�
H����v�.�ѥ�n�]Ux��D^����ї��ox�%��!�����NKx�#��:LۧYf<�0�W�z�4	ռ\agM�*�L��2�^caJˊ�:������Z�&���DS�zu`;%4��P���f�e�`�c�wH}�*6@v;���9_�ġ%�]���gƷF���S�T��0��o����� =^=�
���"�����P8� �ױ+^���#�3*d��T`� A���F�>�o�{�҅W=���ʾ�3�yq�z\�S�Ѩt����):/���G�*����fZ�5q^�3���XRg��X?��p�O����7p*�̄\���-��d[�P	M(�vQ���nS8�Z���j� 4!�f���&N!���[>��^������c���
��Er����ֻ����۠����q�c�]G�1}WUv仓!TE��d�*u��㴧����ag�1�Qz���,���R��yI�u�(֫�^�6_kk���	h<�"��Dk�y���'�ߋ�n�)�k�K�ngX,�h�{�]5Q{�q%��:�Dв��^ndH�P�m�R��
�>lB�D"�tf�����^O3�e�z�stX�g%����u�	��<�W<��m�Y� CDhkX�� ���fß�| An�G
�H��`�h"���L,���;/sC����HL��/�2mnM�� ��G2y�d�of��;���>$�����m=SfM;��&��n;	�,ů�)�Nl�]��3잡�.[;;˦��Ť��Φ=w�^��i^���`�#I������X$���}���L���l��4
��~Ti0�l8 z�Qٚ�(�~�y��H�`i2�>a�S��U.+׸��L��TO��<��u�@����#	�m�s��ӆ�u��*���~��fj�6���>�H+��m�8�B�������l==F���t��'Y����eo���|��$��tT
n���W�k#e��ND�\nB��.�l�,���=K?����p�|[��5��O �x5�L��z�L��Z˹H������ׁ�3�F�Q�Mr���4�4���2k���m)��4e0�$KufN���'W������L��3��̡���i��t��nQ�eJ-�X*\p.22�	`^c�9ν�z,p���ş Ɉn�}# 9|z!D�!J��W+�g(̏���\w��>�����	�O1���.��p���׹��\�h�(6�3��d'�jMk�XC�ݺKc�E���$K8s�1����m0�# �
�Cln�#z��gI@�gAЅ�t���:�g0��Z�2���	�1�6/L��%���I�(.-�}�g�
�)ޔ��}��_���OrV�^���xK(��Fe���^��"6�w9=��1�k�k/s�bQ�1L1ԃ<�)�N������uac?�{kQ���>��
@������R��m+q��j0ߕԓ���	&�Л�軣����b[`�����\�:��s	��G
�� q��H����r4K�;@��]	�D�Ӹ��$�����?�	W.@���)������%Eg��G&�Z�ɫv!%�h~�=p���~xjX��(�߲^0k����W��/	��kмj��P�
ʑ��Sv	�E��1~��R�)+L�
Y�� �P��E������=���WH�zq��{�3:k#� 
<.���?O��H�v���܍�M"r�I�c(��A�5�Ŕ����،�z٣�B5��~��tI��t��X�}�|N7pf���M�ڷ<fțP^�̙\}&�"׏L�p5
x�R�1yQBxV���v�T�%+�������j�n�	��E����#�}�z�-��S��G�=qN���P��76��2y�ɚ�����pQ�XW���4 ȤhS2P��+ZK��s؝ڛ��o�'���g����l~�`�f8)���>��z�����V��������?O��4��o��A�ΐ��&�d������^$�0��ٍ�47.V����9��B��OKH��<*S�����Gy�VJ��Eu8������\����)���kYp�<�l������'��|ݻ�NA~�ֿidC�量s�Tiy�E��r��x�?>W�F����N6a^����}̶Kn��
��-�����>��ݑ�O���ܡ~��3� �(��p85C���pR�n�{D*�Y�`e���zb�1�L���a�Z&�AE|�/Q�%н��]�d'�� �Vx���X����9ݵ/��t���n}"���%c�^�����u#}tD����@OK�IT���͛S�&��#7E�bή��>����գ�$?�o.��Y����DYP1Ёt��#��d �	�F�7�o�vؙ�s�5DZ��[ �w/�E�j�A�y����xR˚���cGe�����rO�I��d���r`�#��7�<Ʀ*Rv-:vE�ُ���?[��N�l�`0��_�����/�����4`0�Rp��3T�z*[�'�L�:��{e�]���z�	��*���I����ފ�j7b��~�_	���8�)��PV�z����D��8����Wdg1|�z� �(�߂]uB�p�:�%��dS8���Q�B?WE9Tt��̀	�ǋ�v��7��,Ö���ip@���ڷ��U�s�}sk���c���;���r�>l ʾ�����K2����"\ف�{>�!3 E���o�.����7��D��vv;��Zu�b�&(��_��eD�>2�H�TA�E#��s�"FhAb@j��%Bm�@�Yz��X��'hN2>��������M]����>�T����.��ʂ�`���<!`B�ju��`5r���`"��$	˔����T�F@�m�\�(k|����;c�XS�D*�}{�!ODC!�x1W`G����a�DG�z��B0�;�]�!� �q�F����?�8K�I��0͠����0�C�0\{�>�'@\�Cȕ��P?z]�*�1���e��C>@2e_���(U$���#S<0N,�t��i�;������'z��'�]�cDm
D��#+R���_Պ�����a^�����J9�
S��%t�p�������9�{�F�N�ǂ��;=�?����_E����g�Z=��;��4�2 ��)��\~����"36�(��C� G�)��T�pN�s��*?O�͂�rd�Л�_&Ϣ�{���vX�v@�;Iϻ�^��tP�����p�?�CG������+�D���o�s~����~ߩ�Y0�4��  Kn	�T ~} T��a��u��J��}Wn���NRVՓ�v��#]��9ʂd]�,Z���̭L Ț ������E��,�/�DM�/}j��HI�O1��س��m����N+?v˶	o�LQ��6�W��@\e�p��uZ2+7�&�����~!OV3�\�Q�c�0۴9����wN]C=��%2�N�b�|��ׂx;����t�E��4L�+��j�d6�YO+n�YUMP���ɜdD�=`` TΙ$(I D�5��^8њR���d�e�ɰ�}v߸п`Q��?��{t�LF�/��k5�Y�#b������&� �iw
:S���\�Q�vQ�a�(��Ͻ.�%�X�z\]��J�K4��}��<�ư*9��isx����?{�㕙* �(��z�׸��Us��:^��]V3�M�߼?�g�皖���rS���jjS�s�g$�e_2'o�G$�����I�w^��'Ӻoh�"��^��W0��rK##��9;y����܅,I� E�ӴMa�sv�!��?�t��� jG�7ښvD��΅�����t����s¼�0�������f�t�7��(}8�"�>�����7��fTP�Y���ٲ����A�T�t�]۪�pq�఑$JF@�@m�M����]��P�7��}���˽S��@O�!�ҵ��n�׹̈́K��X&)G�m?a�S�U#ah%��	��(��+������Gyw4�L7�E�;�r�\1W�}������Rԉ؋����R͚C}Ύ<���:<�����q�\����	�d
+I�~y�<xxQc�F�&	1j�6J¾�8���,r�z�]�U\Уv��.<�M�]���6�����I��B0�a,�[-�����C�o�0�qcè�����t���m��y��`r����l;[��j�7����_�:�����°ԝh��l�k�^;�� c�eIv��9�~}x=a�{R!w&��ݒ��b��v��gO�����\��:ټ�?�[Zڱ�i�	$H����;�\3G�s�k��"h��]3�oz�&@�NV�	B(����s8�WuM���؀zw��(eJ?����,͎ø�o�����1/�ʙNك���A�]>?��bby�H�������OYjŝ�.~M($k*���AD����9.Mn�w��sۭ;��WJ�u3�j�o���� �8]�Z��Ͳ�`�:��� �1H~kȃ���h�g~ã �m{�xJ�}���f�;_^ܽ��<k��>m�&p�h�������1SEi.Jƚ� |N��0� �#�i���_e����{+/"4jS��O;>��g����rAlP������/>àÛ�Rʓ�`��r=����*�U���G4��_fx�"�Ǳ\�X�A�9۱n�5���1��kЎ��y�-��9�1t��&�=�����hN;�}�.~7o�qU�+��照E&�V8W;Ͻ>{PB��ދ�z&'�������	���t���LgO
�,�9?{����@��`�7��������!���[�ʔ��H-20f#!)�99R�4]���IQ�T��f?� �o�3��>�%X0{�}�R�2�GK�W�5�l`o�AK�4H/����dwh�>-�)��o�C��.�r�C�f�����^�b��,9Gc{,^�9���9�u3����o���&�����j������-�T����،�=���t��������`�T����=q�����bff^���@�ԧ�m������_�ܱĂ���H���vr������=�q	7�Rg����_I�/-����|؛�>uɯ��BQ�o����Eþ�e�����A�!�;<�uz*}�wa�N�����&wr��?ȟи^�v��`��ԺP��͂�OB.�,r���	�߲���q��9�?;�Hs1��s��#�U�Ӌ��*��2�o
�n綱� �7g��J�-��u@M�q����"��ׄ�v����Ղ���vW�T�$������S���N�:~k�m��Tr��X?M��nU����a(��̅��o��i@��[����pj�rNpX��W��?�h�2�2-���`�W��/��*����؜Ps
�8 �� @��ݙ_�c���5�FL����;qA>� �k<~�Y屼�G���ōv�Y�7\/䃧�F�J�8O��.�Ҭ�w�;^���ӥ���64_�����
�Ƨ�g�l�N�]9�z�N$Pn�v6 ��ƤK�@���PZ�N����fM�*!��}]��`v����

 �)!���2CJ�����L���Ӭ�>��뭠7���;����@��egXa�3��ay4�w��)��/|)u�4��3��]`c4��<Iٰ|ԩ��T��Z�#�l���q���^�������<r�3{���;"��
Mw�����k���L�j{���i1ڕC�ch�3J6[�#Y�
�o�i�f�u�Z-�@���|�.�g2��L>�	����ʰX������HreA_�pw��[&�����_�{�Wq��pL{��U�w"��RMk����2�zœN<��>�4,M�z�B���~"�_�z|
j�l�T��Q����?{4�����~N�_�ƢE�v��H���ϩ�#��GO��M�/�֑�k�.H�s�>\s5��I�&ڇX�̒��g�0���u]^;��d:�����S�K@�#L�{�od�F�,H���c�\1sZ)5���u}�{B����L�5�?�T#^�:G�-z�u=�ь�FG�C����s�u��j샱�'��|��{���C���|���<$11��];����#Ъ��]4;�V}s|�f#���|НS��� ��m�J(���t55��E��8���K�=�)N&�}���U(�ׯ���w��(����;�%�RWu��J�Ś�I��~��KA��;OV�@�~>���TI9�cz ��*@���򈌴(��	������{��Ps%�n�E��轶g�;*$P��U9��5���_����wU������޲��*�w߬�P�D"��f��"��\v���i��T�ſ�D����'л�?�?�c����������!��*�r��Z۶�+����8�W��N4K����0��P�=A�Id$u�ߪ�-�S�y���m[�aT�����Kw��x_�ȷ��j�������hg����=���������7�0�4�1����@48�Iix��<$���1I��gb`/�V��R�l%��'�H%F���m��=����[��=N�\|��(��	/K���J��γkpۆ��ew���&��r�1�Z2���@`������lbj��/v>��y\m�@�J�0�,!�r*o��)<���QqaaÝ@	r_˦K�d���$�����k��m�=7�8�a��.ľ��S/�F+d�d��]���_���9K�9�ڼ�KO��D��sh�����=}|e[�K9{U��햲>���v���8�O�ʥl�U[�Hx���$��Y�/\��Y�$N����F�	}}P�!���==2�:h~]����y��cQU�ք+�5����LE礮ŭ���
�&3���O�R��u���`HUE����;��:(2S0���1�|�Z�RTW�[8{0M*���+Aj?���!nm�4��&��9���CO�ZF�v���|��.�^�kz=����V�ϰi��=�։R7�|�!hR�� �Ra,�7��&՞Q˺��.��#�vg}����2��B"4C��/�̵4�}�QֻXل��%oj�@�������h'$ЪX:p�¸�wh��	���t�'/e.83}���<.�;���8�U�z�������"���==���ӳ�?Β�:+���=u���oS/������U-���?ǳ{�)9����:}VL5�)���^��.��Y2ri�g1~��em/�{�ȅ }ȉ\�����ޤ����� ]g[�M��޹ժ��q��$�)]����(������)���0��j֧�Q~֟Y����A�yוGEwThe1/�67z�ظ�H�J(�''H��t~Ş*���Ҹ�ϰL�̐���!U��"�Y��f���g -����2���j̞�(�p��0��]���v�z؏X\���̫�=.�jk?��[W�V��o��C})M2_x٘��-����|1�<��JU��''�y����h�P�W�#��������bvM��e�����ְ��2~��N� ��M��F��ͩt����ʼ���F���U��y�\Xp	�Q��uչ�0Z�*�nԔ��;�!�k_��CN��x�E����PM���<��i�AՓ�"
����E����������^��7-�e��ƙd9ʇ*��x��JcJs�>�ԕ��M=�EC?x�#\I�g��3U�{7&��f=�Vwh� �l\l�h��t��+��
8��l�e��h&���7�<���)�'�Kf	����ːDz�r-m�C*d�dl�ou���"(�bV��_���d�#��a�4�`��O��%�lӑ�:
)����X�B*���������RN��
��sƁ��� x�)�+�����.G;�G���q�_����F�(���G�~��>�~_&�6��0`��(�[�\�N݂]\����t�?����s7^���//��s2�PK3��� ����C�FC���K+]�)��GCi�H��tG
���&O�ݕ�bֽ�:^��6�R����$�Ԇ�Ig�g���Q�ˣ�j�W�OX��W<�����DX|�����Uu���qu�	k�Je�Xpӕ9��)�d8
�Q�a�9"=g&���A4��wL�|���g!W�<�fJ����oh@|��|��N�`w�;{�>�r-W��nN�	�M"�}i67���#Uvß���+����eI�~�]�3}�eC �ؤ�qc5�
Z�:�z@��5(.�Ƥ}k�Zs����J�?1�7k����<�����xf�	����^���$U��.�Ս�7���7��q�gV�g����t��Mgߛz���j����Q�?:��������;l���0�l)�J@�@X��'��jwx��پ1`��p����~|�<�	>R-��鞬G�M$�_x�i휱g�i�
�7$ cE��ɸ~�O�T�L�I���o_����´�nI�y�/$J�L��ȆA����2�׿�F�GF�=�I	��a�_r˟ ��P��j��3��q�iL�N�����$��/r�J�o|���~��bMuuC��E���%�[�*R�{�����ĭ����c���όI����K ����u:�45��i㫴x���CM����8V/�,1 F(sa����j}W�I�{ZH@ڃ�NL��zxA'9��p���PJ���`|ĩ�֒�h���CO����t
ujL��Y�7�a����6�����w�o�x�3R��J;���t��h E׸���z���7�KX'�x��ڢ�ULW������ipw���x�M����^]��;:E1�b3�6��t�'�OB[�0B_�i�6���,���Y.L��y�ܙ�F�ouZw��O,3$m�r�}��6�>Cx#��t��8�����QM/_ߨ�c��X�
�DzWi
�;��^#��HWz�{�� ��.%AZ(!�����9�G|����u׻�k=�יٳg�ޟ�e&|gB�/�!�>��	[�^l�I��۔��<$� ��rŒǅx
-V�-��T����T��h9�	��oXi�&��I"���yEH�;~�.k��b��MԊ.l��d���u]���m
��3�����8'	�Z�s^eh�����<9�hW�!j�S�w+GǪm����o���%��#*��x�������i�]Sr�ytfh<Y]�4��i?O�R�/h�7�$]��ث�f��\W�=?.-3Z�X��e�.5���'��8�o���7�zj�3_��g�E-S�a:k;�o�3]�Q�j�����������&�y�b�kJ�:%�h�R>��9�!j�+���� r�)��(�8}�S�۸np	�}-�hI� RT�L� ���<���fH��n����``դ�+�r��E1l<��
B���LrB����G��X�c�[Hd��<6�� �/o�M�R7.u�����qt�i��ǰs�3��\��h�#��ʇ�]�k��|~;�L��y`�0'�D#�L��J�""*��#r��6)�^!k
�����`O�Y�0�m�[����Z	>'�g���])7)I��\��6��*��8jO�SjB�6�ȨUW�m���Z�=��6-g��X4OK��K!i��@mx��=��:@����"r��CE��"��i23n��FƬH�S�U�Ca���m���Nc9R�i��,2�Rk�4>�y&���H��^�OR��cl;���*Z
��Y���\��&7�X�s�@��w���Yw�~ W�Wǵ:���E�B2�s������m��#��jz�}���rV)�|+I�յ�y� ���7&06�5}O�U��/�a�+�~�b�m_ �f'(��޵_i�OR\n�@`K��p����>�ACf�d�<�j�wgC�_���B�)��6�ͯ�ne N��_�FA�sRG�{ô��� >Qį����U��:s�zOp����551y����8́�����G�������.�k�5o&���(�Ɖ&dd���F+�q�=�Y�"L_�G"2,�T�嚡�'��ܵ���)p�`��p*o�C�EB|s>>���!}t�挿����qZ �\���mK�W�G)��|s�Ɨ����s��k��s_���d��#�B7�1�
lBR�EH�u
�|���ǝ�Qe���%�Ñ�u���J��%͸�4��O������~�"�͢����#0�OHK�ǃā�8�ǀ^�B!}S��F����Ȭ݈��j�ykG{�A�P㞣x
�o�USu�Q�[��ټ��!�
e�T7f�<bM�īvk��ZȦ׀�Ɇ�j�$2��N��&��ϛTCۻ��o�&�k/���u6���[,���6!�2BjK���x@�轅+�,;�2ʻ�n���úL��ب���:O�Yq���5��+]}�0�b>M�[��V5*VRɄ/���ARՈ��o	��<�v:|���`ϰ^Z�ƹ�I�C���ܝ�:�TY�$t�Qr)��}�jM��CTS�k���v�1�諸�[�b��nv�;VQ�resK]�\n�dG����'p�b�V�L����k��m��_���[n]4Wh�gGi8�"RW�h�n�ʷ�!���Ş�$�3�n�w�-��"'��4��o�	�YWB�H��#�3h�D��_�mA.���9̳%��q�Cb���{����Xrz<B��f!��E��[+tX�z�(P�rZ�`��z��*68���E�m�NY&����n��<a}�(�j��Od]KA�vN�>�e���+]�
s���'*vP+�>	�-�6
�[d[��Yj��oh�*�кT�:z;�38߲� ���ƒ�8k�vW�7g��[�7B%�c-���M�M,�*�q�L��.$��$�w�?���=a�Q���5)�$�
ۋҰڞ�}��s���lU���^Dg)Ќt�q���[��������)�&�>��K���6��FrY�`{|QU����=�20
 �*6>��$�O0=�U�Mbّ��L1%ios�<p��l���ot6�m���oI��V3b�xҠ���W��Ob����A未c�[��zq��8$�����:Ӭ��\�o��Bܠ�z'|���I��zẶ��[��5D�k��+��
�J�'W4�����yߚjYE�l�%6΂��{#��+�_#�{�?�9���X ��}�U���n>g��͕�x��C���Z�~�9��ۮ������DX;h7��wH���~�@@��d:t���@��%�P���i�Z�HLLY<su����u	�⮦1���}qa<o�x�9�e�?n_�|�RQ�
�gT�>�g9z����j)@m�T�V�]�l/&�~�r.�*�A�{#w�dլ|�:D��+��T\}!��³���#j��� `��:�$k�ڎ��>0$�<@s�[�9}q
�K5M��$�y���"�'�k�Z���E��M��|c��:��+w�e�@�a|�;l���V擖�:]X�b>TVw/�2{��)��5ta��U����.�k�3��w<���ٓ�ҜD�1$��σVk���k����-�{������#h��6�ŝ��LqVuSU�`kN{�嚰_�M�.��}�@}��ul���Li�S��g���5]�+�-��`YTu��x2.��e�̐hY2�~�=�j(���UU-�7�&|����Z�"[�%���dt��W%Me$��ɒg>|��U}Q���h��{�=�4G_��x%�1�w�^��R�Wy�[�̩h�h��B�[�B�U�r���Dҝ͞��V��-0"(vߍ��X|�����*���*�l�DS���d��Ed�L�[�~G;�f�Z-�ж�%�Ȁ�|�>�~�@��Lh彈��6z��Ͻ&	e��J� LOot�:x��Zg�Ϟ#��(#���.�Y�L[� kC�ի�.������|�륟���a5m^�:V��Q�T�c. ���X�	�BϹȂ�fe����99
/���YZ�h�c���Щ��A�ac�fӢ���ojA�_�b͏��������ߞ_ ��z��I���:/ r}�,��C "l!w,d�{q|��Ǟ�������sVα�m>�Z�D[�N�85�
�m<Q����)w�������C^EnQ�S�w2��X�D+��J��0�Ub� ���Ė�S��r!-f�X:m|×/��R9���7ƽ�4u���]�&�/i���Ѵ�>�`�rX��,�,����q�ߏ�����jk�4�������$S�t�Œ�����o@$�q-��L�`6�L��Aig���gc�ᶂ��p9f���:�����F�i��}|�.��E��+�ɴ��[}�!�377!V�W��v� ����(���fūj1��i!S��w�x�=x<)���!5����~U���)Db�[f�:S�i�4�+Ͱep[5MS-[f;�/-�4�S�mX�g���e�8��E�nIV�߶��<�IR�D�+��s�
H��ZU0���Q�㙹��%*�D�r����-���G���w�����׊h����a��-R�U ^z/�_-�]y�e�8;�M���+_S7B�4�
���Ro�y�m�+?	����\�ݫD*�_��&���NI)�;t��&yñ][+�"թ�!y��˙�z�Ֆ$YC���0�e��[|ح1ʽ�y��OM�zܭ��|q����VΦ{U�Ѻ�z��֘��XS��y�"|��;�i�x c&3�ڷ��k �Oi��[ׯ�6�m3=?�U4�ݴu��x��#1�x()=ׅ7��'��B� ���Y��idr`�X�oH����5�2��=K�hla�h�l��MY�^��$�N������Y����*�� �R+����-;��ؕ����kƱ��[9���{o�XV(����P0O~����NV c����r��S�E��"�6���@����w��Z݁�#"]�b���)�(RazG-�UC��gp]�9%�dw�r^)6tt��pҷ� �7��uX��g)k�5��q�x��G�
���6����^K���x��0�c�sQ�&�H����a'�7{R;���l?��X/����
Q�^*ik�����8a^s<e�" ��N��-�9�t��u��!P-�����'�CAէ�W&�r�+��f��]�߇%&a�k>���>֯�����JW���U��Io�� ��^�������޺�ni�o��t�_T�u7-����C�$�H�l�7w`�k����Q0 S�[�f��~��I�\��Q��'�6���L[͕6eE���*�#��	Q���3�R?ې�Q��"4[�3����ʘ�Z���eM"��\����.�4�\E��s;Q�i~�%X��X��@�G��?�9e#�~ �N�DV����X��&;a���L�)��6� b���w�9�����:��>z��w��7���C�5�&_@�	iI۪�|���F=��lG�2R޾�wyJˑ�{{�̱O�_U�S$z�3�O�qЫ���{���E*#1�x���P$G����GƄ� 5�M�'�<��|����9�SLf)�Dn.@K�׬�D7o�Љ_��6`6�^w Չ�� �2�+� �D4��(�^�m������@�᯼E�'��C�șq��d�Ze����D��]�.�+����:�t��ʐ�5�>�M�w;+'v�pX�<9O�������r-nst�o�Ho�P�����ֿ�<�H�LW��Z�eN2��4���O����ؕ?�{?�id���;�9t5|�0��M����'!�O~���ᰣ�	����E�>����)c
KV�z=��v�cv4Qm�]�%l{_�/���J�z�DԲ%�������T:�G�� ǂ��-�k�=p
�h*_.cr)���b���n��B�����M����ŝ�@7wT�
�*�u}��ļ�>�Hnd�m-��t�S˔`��mX���?'[ǭA�64�3Q�E��u8Έ~t5xխk-h�3��	���f>�9�r��i���t�m�W��x(��;N��&���C�ig�L�K�yeMHJ�7+<��T�I�������U���o�,���[U���@l{�zh_+��~��y\T{�Z|
AA��S$:w��	!�YUa�|�u��C�^U�Ms�����Z�Pqc9c��V�/�a)�
�~�F<|'�6%�jk�)��@��v��x����6�E��EK��+�rx��u|PH�	Qq򉶵�{�T����O�ԽOڵ\pL�Ś�%��S}��pKqE����'	U��8VP�s0��\:�T��5�(<��'�K�Ι���5.�������"��U\��H��"N>X2��f�p
[�e9� OF��4�(ܴ��ͼ���)��t2a���(��R]��*�
�2y B�0�,�
�I/�{_/��bsw�y���??~�U[a%�3`+��կ�DU��ǧ����>��1Q\��
�l�����<#u桅'�G��3�������@��:�[��Q���a��N��м}�Ĺ�*���&W,���.�8Җ|�t����%U�Bk;ij��gpM�̅�v!)�\o�g*���bm#I����a������P�!;�X��Qvn3OU�L<;���tENe�[�@fv�p �%��s=yd��ѥ�~��]�]ҹ��N��k<YZ��Tl��c1���1e���\@YL�Pop�R �[� *�솆C�XS"��R�O'� +?/��$���U����N�z詡����-�Ƀ�-������y�z ��`o w�ne����~s�>���2��Д����R��+K�M��]��tų�Ӽ�%(ķ,a���5)n>5ޣˡM���	>��4���;��N���R���2��R��&�b`�\� r,s�����e�$��D2�ɑ���jUG���{i���XOmu��[���T܋�3V��%_ҝJ^�:K�2�����ƻٳ�P;\�~ϔG�)�Н �|���R�����m��r��[W꼟�Fi���ɯ�6�|�^�^ee�Ʈ�trL~'�݀���ee؉)e%�X�����u{}N��:�!��l�4��n�c���b�܉m�?��CN֖̂Qq�?��@�^>�f�&�ȃ�[o��M�B��M�"xj�O���l�=�������ǣո��x
�iǩ8��|��s���׶8iw��L|_u\�����c�"��il�1�>?�*5O6O�@�����H%r��M|P�6n;o���-8�BK%_	I=~܋�ۂ@HSVAeU�LV�򛊷�y��t���=ҫ� ;_p^y�T)|Y-ϻ����\4!>��z�B.�|��҅�<3{z��Psv��Y[�Ϗ� �L�6b'b��:ې�싮�,����=���7�$��,'�1w$ׅ����C��6
@�9�J���F%Bt]u�*�+���4�#@��߿t��*0�iZ��!a��I�VjOc�т�qq�K|9��'�Q.4Wڐp�~���D��9�I�)�y��N�
Iic��  �A!��n I�p�`�p��[q��9���6�HV��`�WF|	AVMw��/��H� �QTJ@�˶+�Zt��5�f׾�y����8	;`��H|���a�zk����'ʧ처�S�v �Z?fIﭠ�1��k� �X!��e����^c(D����ߊ�y�E�A������F���)%*J�H~DR����K�I�,ѢU��A��;a���j�]��-� �0��6�%���YEb=xk��5�Bt�h�$��R C9���N�����ҧ���&Egc�)��7�:�(uaU/(=�H)<�ꂊl�\^����L�D��JS�G*!��Թ����6�U��O63T�����R�W��NIt�z�sڱk�`0�-3	 N�1y�S����3�"�꽡Bg�B><4�d{�$	+b�Xez���zԞ$@�	K��2���9�:\d^_�݃"�u,Օ��n�UV��Rd9��s`6w9[�� g�?l���R��c� �h���cB�b�������^��*�q��9N���*vLZ�������e"	�أ��Kޱ��$Ia*g%��.��9���mXj���/�1�j��@p��d�f񑈂�dʗ�X�S:�l�.f�w�e�u2�߾�dr�}�<(��1���k�}��sJ�Xm�̩J�.��`�GGr�ԉ��@����]3��������^LG�e��O�2G�n�"�� �7��aʬ�ry��7�ۼ��}b!�����Ĕ��e7�WW�Uq{�H9)�ޤ����O�b�G�x�T-�gK�'Bh%j�2��>i�����ȴ�cJ�/De0[3���c���p��'����ȳ�N��&���%H�o���3s�u4)9}|�=�*�,qV����߲{�+�[���_�L��XGY����d�m�nz�ƽ��%U��2�Yʹ���c%$��Y"������C�=�`���Hy��*�C���@���s*R��CDÉ���Д4��� ��9|�)��׿'I�.���/�g�}1���������,����j������ ������~������I����w^b�����^����?#���S�Bw`�������86�L�C���0����^���%���|q���9=d�4�+�ލ�l��!��]�dϮ�Y��5�:���-����%@@f[�J��'����@`�Z4o�k8gԋO��>�F��$_Uy��D����L���o�soߤ)Qˍ�1k�T*���Qd~����'��<����c&%>�:�=*�k�-�2[V�z�>�f^���4}'Xh%�3���Ĺg�X��~�~0J��d���po޶�ŉF&)�CZ�&�'H��JP}�<��f�*'ihV�����w���D�2����}����C�AA���Z��U���{�3��߭2f_�N����7P#:\�`�[�Z�ïa�8�}�+� ڟ�*��Y?���pMv_)��2�Gz5Ri6��t���:v1^�^D��lk��Z��$Iվ�WJ�܌�v^K��%li����~\�x㓈�v���(�!�8���w;�E�&�T�������
����Z�+���^��s�c�z�A�Zk���[UM{�����{�a~U}	�g�0|���RH��^��� A�|$�x�*�Aά�����"vW�n}#��r$Q����@v�&�4�[{���Y�غL����M`���Q$�|xq�xR���#l��#J6nf���̪�J����7�V��g{"���@��}�-|*�&	��|�y��
8����s6�����e2%��
����X��C��}�U{�T��
khO��
1���C����9�p��
^����:ع4O(�mJ�A��g���!���{���+�M3��fP�w�&�OG?�|E{Y(B5\m�l[��'��l����Zo�ը��
�����aJâ��K�M&5�-,��H���md���<�j||>"�>_�T�r����~Iq����[�}��Hy�(TM&�`��i��rGn�t����,/2R��!c�V���{��{��۲N�ǈ�@6p��&���z�F߷ �=���!i������S�c�2!��C�%Ȃ��;z�b��c@6X�=�j�ve8����4i�2sF�೩����(��"C�À����a���`�����pn�NV�H�p��C�FDD�33Ծ���h��AO��+��e�&���ѓ�)��|ȉ�B�rOxC?��D�����9@��햎ײ6��c'��y(9�a�v�hV�黎�X4d�j�;�����+�v�T�����8�#Q��d<���õ���-��C��&���cD\D��O2�����+�`��J�VP@�́��Z��!��6�juu���>-GkX.&ᙑ��0�hw�¼TRp��W �W���u{
,>MaB$i�R;2rr�Za岦HUϖ� 6r���-Y�tH�;+�e!�������wH�@��P��|V#kV�ݬrO&1���8�ٺ�Iص��$���?���o�lg�I��D>d"���L����hM�b�(˚{
���ha�\Z4\{�*4�@n����k��i�o.���8	[�t<��q�(C�6"��T[$��$�d�~6<��RL�(��Ob��)��\ �J�]CB9��e���n��,��4Rqp�b����gٿ���T�=C���i��{�l	�Qv?��Ņ�W��r_�C5��;�K��V4���0�ј�[�﷏�=�[�٪�����ǻ�Ʋ�~=y�]�9-]ћ��f��f�i�̺!�	�b�E�����(w햾�w�Oy�_iٵjﾹ;)���}|��8jt�Qvɦ-� �����OD�����gt�m���'�䞻����!'ݭ��ok���W��Z�N��}k�L|k6' ϻ��~�����銿P?v<j�J����?k��vtH���J��x��*D���E��.r_+^�����D���+���$��[f�;SvW����J����t���5�����U.j�	' �nw"6�@�����0�W���,�+>
2��씎E������	���QI���0��>�ik�N,��U#���p��r�p�ũ�V�}����o�������� 'q����,����6�kLW'rx��e�>'Q�u��j�����S֛��������a �7��
�t�Y#>��#�5}Oj!غ����ݨ*�*%8�U@Yp�έ�njg�ԝW���a�q1QG{/�-0'D��������/�������L�/�V7=^�{:��R����v�cJ�h|���\G�,���SSo��*��Y���d}���iX����wT��&�0��M����� ��U���jq�6eA�����|�H���B����� ������!<.���@\�j-$��%�^�9�M᫴/T ���ơ��;�}Z�Eҋ�V�9Mm��և��ߤ������TdDT����i�0��9�(�U���YH\p�f�ïL�<��,�����NU�1�bg�>�!�7�W��8~[��!҅���<o����}O��А�]�������i'����:=2��m�^�=�E���4;��z=W����t}���B��#��%Mb+��k|ޡ���	��@�PuZ�l�ע+Wv�y\�eWf0���:u�i��b*p�}={|2$ry�2_�ʊ��7���5��1��&�ۯ�����uK;���|5�=y��4�5x�B��]T��y�(B~TOA8��6���$N�p�ˬj@ZyvHh��jrM(b���i�>����(���-kr�TŖ�����u��Ğ��*��z}��k�6� ]	K�~Ř��p������=�.O(��~�[��Z�����\Ӣ/́��/�ii��yը����O��%�[A?�H�>��䞿N�%�8&�IW��ү~m�Sǁ/���ܤz��qG�Y�,Y�n��ք�zD�!�����e>+P��vʫ�~�=������T_�e�>��|�wJ�"��z`�T�+�;Ojգk<ޱ&�]o�Ђ싮&Z�2Y����D���)j6��p,*��֏�|(�@���E�?��M_�[ �*\����缋��zE
N6���s)1��6J�6�������rDG,���x��Y�Jջ��iЂ��B�|n�E����2��4,�iN�Ep�݌ii���T1҅T`���]���W *����oUS����ʆ`��<X����3 Xx�b�@�!�7�\����!�!�4��3T��hF�Չ�bx��M�}���i�K��+��
���<i⦛I6NCwz��m�v�F#�R�r��5����y}ҥ���7��N`�*��½���s�O���3Z{7+-��8��ֆ�V��Y��7<�i^��;�4eP�a�hi2�2���ᕧ���~J���<O��%�Q����%M`�ƣ'��9c��)�.Þ��Z�*NÞӒ���g�6D��z殍�:;b3�ӊ������n�e�秫����\N�`�9��������<v7���Ƈ�$~o�y���ޢ�:�0g�y�%0�w�Ea��9�^伛��a,�M���;���P�T�)�3l�%���q�>�S�߽ݱ�������]��'�?�)�g26�7���`���D<+.��ۏ�?��L����)���DN3�����79��<�ʜ��%�pjʤuֵ����	=�n}����M�S>�O5'���k�1v�[Ke�vkS�.�����ݺ�)(,l�1�����h�5',q\�MgX!U@�Ĭ���5(��{m���W����9uSS�A��������k�r	X���A>�<+�U@��tБ��=���̵Y�WB[͛�$<K����EL?ui]̺Ӝr-f����w|��*��>W'V5?>%��c�F����LR�u��4ۍTa;Af���G���*��n:�R¹/�|���8������[`u��$�-���,�������ӞZ�0_���� �RH����sԲ<�<���GaR@��y��+	�Wn�?�ʜ����%h�!��(�l.O~��Z��=�*�DI�]:�S�G�`���Nd��������kVb�&gm� ����'Y=�hO{Ƽ��}���N�X���
�����[�\�����?t}�V�M�0C���o�\'�>�P�?��d�Qʨ����1�y�[�)G���j�n��8jf���z&�Q�ityr#�Ϯ;@��IׇV���\�|ˉ
�|!�$"BWɱ.׆(Y�Y;+/�x������^���z2�U9�V;��m͸ں���Z��+�Y��8��>��-T\^��T��Џ�䝒cq��R��m�\�/�5a[]��m,lEJ��Y�Э�4�9�ǲ���c(����_Y��[�d����B�}v{�x�f��?���Q�������r��FW����䙩��r��`8�礭��kK
=��t'x���-�p���Q'</�+))Io��N���O�b��A/]����j'l>�^s����Jٔ�hy�ONӽ�g����ya�f��A�C����'<�.�� �Eq茈���O�/ӎ���%i���63�����e�c�~}o�>ͩ__���i&F<���W��i�;��ӽ��J�u}�6��Ox�衉L�n}���>Gu��(g�ޝ��[�O�D73�jڇ�����?��L9l`N�~���@�J���Ldtt�#�^)��� ���`ϵ��G����՘A�{~�]i����z{��3ix�U<1ES#{Ү��Օz�E�i$G�׉j��5��ΏlG��� ���QZ���B�]�Q}�~��Դ]4bc��X�s�����JK)X�y�ݑ4ϬfEۈh���Z� k�iJ0��6+J�~��I9�3�1����)������E��(�ds!F���pv�쌘5���^���y˹��4V@��f�b��#\�~mmm�di.��$E��/��;i~dH�'���kЍ�&��K`0��Ȅ��$v`T9������iJ�w���]nz��?�9�iv}�c_D#�#��� �:�����N�>���L��c8���Xdd�ܑe>�<k���MrV������P�;�݇�9z��`�Vs�P*�ƳcQ��=;;޾�5�y�.�;9bؔs�ڵkĦ)^>>#E£iJ���-����BQ)�T��Shcy����]�X�&L8��M����P�@�k�#��������QUMmֳ�d컿�q�<1������5S_jSߍ�_���@��5���1��!�6+�MS^�!�V����f�L$f�/uf��)�n�a��]�_`5ݹ��3�4P���:&s��۞$�#�7;e��t�5��\���gmy5�5k��$Tf"�C�'ݺ/�w�^\�|j����K��5-�*R�@�7ä#n,J�����p�NJ��� (l �!�TU	w�^7�t�KH`��l�%9��_?;#�+ ?6��N��g�Nv����u4����e�d ����uj#t�jCG�l
]hQ�A��陘�\io>0�244�Ƹ�O����t��ׇ�\�Ħ53X���1���dB��8c�O3��,�ç M���K�����0B@�!��R�GA��۪|Ǧ�� ��T��$�۲�w�G&� @Q�m�!D��N�.�y�Λv:���`0M۵��ݑ������@+��6�e�7f�SRRz�R�(�Gp���L䔖���!��e���?��F������FH<�i�|�y��n�%�,/�.�y��1C�-kdj�/x�HR�ABH+q2�;��}]A�f��<�:_���jW�/s 	hӯ�B߾���<ӛ,�ׇ?و>�ݞ@�_E�n���^�1����E4탊t
�O9�`�m�h4xm0n��]q�{�`聑��z穆`��mf8X��w����!t�;ݦk�w5�1?7�K��������"�[�SJuL���#�c4f��C���0W@� u��y�ޞ��Q~%�X9�!�~��+°�gv�k8T��y��<�"�i��xe��z����i~��>)""bfq�������ג$���`������?��������Z�ciP�a�-jj��s����Hg�b�e�8��4�d�FW��ו��Wk
��.N֗���</�{7���B��<�#[��wt���r�4�Hp�~oy��Yb��)\s Ja����a�!��K'�!�F!��ԿkN5��5��f9�~���fW�A�B����;�q��4��#���5�%��y�ɺ���ݼۍ������,.l��m����Gwc.ǜ�>J|� ����̧O�0U=����NN �0ź��Ͱ�wu��n��������i�����\j�+�9?���ܻ��.o�P�>|k��33\�~��S#kQ#���ܝ����@��XǫS��aL�!��g�ai��U4B�	��e�c>l�1|I�N�X����7�1}!�ߩ��s�{�������xえ��ʭ@w��&��-H�w����[I���΁?����.��~���j~9�k�_�\/�:�Fs Q�#{l���3���.����us��=dJ���J��á��GVN�WjD����"��O�?ן
=�ރ�0�a(P
Ŭ�f4�72u��F��4�,s6oJ�(�j�� G\�%աV$5�cI�'�;�� �#��A��i1�[_Hc��G�N�`6�N�W�68���!�� [�q[��Ą[� U0���s�Y﮻3��̑�3^ 7X8�:|bpp0P��� `�����fA̛f��/.��{_G�����:��*ۀRpv������	O/��A"1t�]��JO�ز]��׵�k#�#]�ă��*�@f��� �6�0��U�u�FĕK���~7����y��0`��r�գ�-��uu�&N���l�T���B����>bȄ;����*�s7���s�K-�#�K}H���V3E�B�w�q2�1��o�\��^�4:qFu�R�̐V��iAd2���%�.|p���S��[�}����AT��Lp�]�#!��5*��pM��Xp����#�rt�$���Z5~��>�	w�e���C�B>�(y�i���|�ږ�C��ߵ?y��[�D�`�(5�"��i;ފ��̯�@j6��i��V
��_鵌�Z�o�d�{W�<~���E�#h�l��$�\jTS�8ɥ���Lpв/����s�QGBنPQ�EA��7!�����k�ZD�+B-�f�c`޸��t�"o�T����'T#8>�F�
����W8S�����([U�F 8J������k<�o'�n`�����3��kߍV4B�Y鎬��ݻ�o��A��7��N�T-�F6���g��PB.;�*��J9�+r�/��yF����X��8���zn�T���G<�QA�a���ܩ�a��^��,��
v��/��sFiՇH���s��>�q�'+l�J|�1�d������B�xvv�DyVPa�R�e�0���6m���M]<uȱ4J�c���X���ɽ�eUs�dnGAv����p�� �R����9E��z����fEw�W�@��.�1� !6I��b!�HH�R����5.h��K�0;���1�wO�"À0����N�s&�1��5�F]�Y��Ai,�Xƨ���2�ʉZd�&F;{^���}iuv�{s�3Fri�?r0rf��$H[�0ȌX�D+O�;�B{��#�6[3�x����V:�@�Vz� ��:��X0�r��2��'��
˄*{Њf�x��	O�gb�N���O�t���7^~f��B�|���l��o����D�*�R����l��/�gEWk$��r� t�OL��˭�9����i�w\jN�\ҫPS�4�*��6y�`��CM?ɛi,B%$� ��j���oȥf�@���x3���#�;�Ԝ0�A-�.A'#f�VWW�b+���m& pU)�rt���f�I5�yp�<@r����� P�O[m�un�D��v����$�Ù����v�����*�I���f- H��v�Gieq�(�xfZ�8��ˠE��w?�a��0�������/�������C������xV���X���R)oeH�D���>�7�D�ĿI �f�������B�P�_��kte����
(��M ˰���#<ѵO���Ȉ)
~ix��7�]�]��a=�p��������ֶ8�wx��r���QGy���/S��	eh���TR�_���,��@��@�u��31a��~Y}���'p�w�^�����`C3ޕ�~gL�swt�%5�H3gۦ"��2����܎G��.�|��?�.��`�/�A,I[�z�4��eʯ1�+�s����8WY�Ɵ���IE������	�i��+�R��p�6y���N�Ǌ97�Šo9����!<I4bsrA��+h]k:
��5K��J�L�S����:�y|�PF���O?�mɓ�X����_�'���yY�/�mG*� ���$�d�T�p��d4��?(�%�nx,��)�+)� �o�G��d�F�E����;��[�*#���s�L�~.�%���lu}eBr3�>�t�n�h�z�pt��Ȧb�vK8N�`�2<��F��3���eƺK�d�te����6?�س����{�G�7��e i��x�r��椄��Q��$(��P�}>IS���%�'����� 	A��Ί'R�q��3G�`϶5N�bHT"�	��PWJ��A�/�RM��G����EN������
ZX�X�^�i�_ڒ��`�s�\U� ��Dg����B���3�&��&�0�+c�v��\BQ�v�`|���Y3�_�4�ܴ:�s��]��/��iǀ���|^瀚���)p3�!����_�T����_��_2Pל��z�+��?A�_�����s���1j@��?~�e}!j�B�GG��$��?Ww�O���i����E:������6}�:�ԔRO�޺����ڰY$Q�8W͘)���J;s��٢��SCr��z�h*G��@��������V����{q�j�.,��ڤ��࠺G*�j���[�>��ͭ,�V��&#��C����)�;Cھ�OteJ[���D�C�#�#I�LD~����������w���Sh���ƛ���d]kh��
�׈���F�֫�5:?���&�4���&�E�ѕ���W�]1g�hҢ���}�-�(3�#�kلL��`H�U�ss$��yh6�j��[J�~ֵ	9V�[���f�O�'�O��K���eX��Z.��ҒJn�_ɤ��aF�8C��M��@��4� �n���7��}]�]����$4S;h����Eú��]�5��_JF+�90��r�:r�͚:���s�Ṕ�T���
�l�j��}v2�ݻK����\3 9"4�u�ɝ�\:E~s$Ƨ�}P�>��K]�������2�,�+̻�a�S�ow�rG$O[^q��_0�t�|��k��ނ���'1w�'�row��H:�f{M�U:W�ƅ�"'w�;H�֜���7vp�mR�S%bg�y���J�;�rJ�y�'��6&�]�:�{�ѧi��{D��azU�Z �yb�ۃ�:����'C�[�8~ћv�Unx�Nϣ۠c��_w��s�=/��r
7���gs.����PMfQ��#��)�FP�)�;
�(D��4�HE�A:""-(ꠔP(]�H'�z �$�������]�w_����Y�q��s�>���v���\lUu��n����p�e��^�i�kWJn�b��4-��/z:����{�y���hK���q&�j��|�{G����e@5���mR���ni�q"n?~pb+��cV
4��� ���58�w�����Tg�ON�-@nn�Ȕpt�hB2�>Ι��^�m�c:���f��n�x kr��6��M��{��n.���]��	�^��;����w4������(����?�D��O�?�D��O����Q,w�}��t��������G*�a�j��8��ess3������.S>�.�6��E �M5;ח�fw��<G}����
,�KD�r�䕏(V�M]wi:��Qz˽�w�ƈ[��N�}�<��HS��ȃ$�Ra����
@:e�I.����x���pj��E.����͔p�4(ES,w�5>5S���_��Q��թ.��:�q�d����*�]�O��_���(��.��k��B=�!���|U��5B(��t�X���n9,�U�P�0��f�O���Fn��g�WW%����{��}n����W¹��~��O�
K�����=>����V^<�${�n�۷o��~5�T�P��RI-��um���dP��k��9c�4qM�;y��^H�/^��@��gyp��2��Í�Ύ��ן����.���<��}a��dT�_�)/]�F�r��)D��oom�ඬBH��<QUES ��HҾ���k �=��q����;Z��j�[m�;F�����	e�=��%-�g��V@yG��*�_�П"���'��FH	���\�t�α�[�Ł�2���<K���w���~���'kO�	��Úl�p������Y{T��2tJ���H������\$!g�7v���1�����#�#45��^��@�!�j�5ߏ�Z��A��0z�֤�hȔ`��LW����`���!Ͽ�0O��No0�65���]L��X�ʽ�&?���ի��mi�j�,� ޣ���D�%ni�H�!��r�cD�`4)A�љ�<��n�����3�a7l��(pUY��u�8��"qi9��bBi;m���IF֖�J�?�)�:�G�G�r ��sjϏ.�˯΅���\��2A�i� �咱��&�=����DG���1��_�V�yɸh�;�<D�x��y����It�����0�#��xM,_D�*t)�f�K7op}�%�q���a����m:6|
��1
����
�?z��Z���!G��l�y��,��b+><q���@\}D /}��~4���1:\ӟ�}��h��?rZ)��u��4g�����u)Z_M�zN��; �E~>-qͪ0�>u^X�M�M���Z�l�%&�ż^[��lME�Ѫ��PNvRMJ#�F*[ :#'Kp�?��yq���l��g���$4�1�fu̪��*������N����T�ՠ�'�k���u2�د����[#����jl6��p��+���u�ܕ�A��Q��oȺ���E��L�����?o��JQ�BQ�ZG�
�[�UK�]S��#2���H�����x<�.�8�5d]��{���
�zN
�覻o�����\*0pjE�}�@v��}c R?W��w-�p��v��8pbǥ�};�����������_��y�����/�<k��!��`-���Y�l��dԗT�������{�\�דN׾���6Ɂ����YJ�vk?>HG��sg �0yQn��k�4F$�5Į�b�Gx��U u$H�>�]�k��`�<�c�b/o�D]�^�����7f���������1?(|�:�N2����1��wא��{'جn4��>R�:��#�<f���L*|ϒ5�x@V��Q�k/%4�
�
�uF���'�$��n��A缢zE$T���������f�\C|���P�Θ��#��RY��819���I�<���o��C�XǼAZh��+���Lq��M#,�X�8N� �4p&N}}������-�m��c��+X{A�������>�=�F-����kLh3��X!�����m{�p�{jf���c�����y�BE�f�#E\L�L����+K-Ǝ,< {n�0�Cz;��\y�L����M��2�����:����Ck��}N����������TmJ��h����u�W6���߻܈���1��E{qa��X�z�*35�	 � ��C���}��E�jʜ7�z�LhC"���kGN?�x�&'��+�C��ܷq�/`���
�������y�J�W�@��EB�_�#�&S�����?����
�1F����ӉK����"�&8�S�[uB�b
�T�2C]+�I��ty����,��@�x,@̺��7.5v�/��>* �/%.�>�V�^w�J�#�x)�����S%[|�/��;�o~� ?.�,��&>|�l3��t���Y��������w*�=E���� #��sI�ƽ��FD)9�k�B:���IS�ݻB�]C�W6��;�_����x��r��y+�I�0���ɩ���o���|Ȑ�F�]��
գp,��Yn�u2r�ע�à����K����z��R�,�tEҾ)����{��؍���6�X� �G�G1um%$L��I�j����e�0�X[Kv~�>��w:p�z���ar���p=�L2:��ݶ�풏X�d�q���]�#*\.�#�ݪ�+_+�2�30�r�j�������<G.�~���
oBյ�]+Ei�׶2:�z�!y�P�����k��]���t�A�TI�����\)o�{@\�F~����2��_�k�^%��(v�_�n|�-O���H�Mhs�z��Iv��}q�k ���mÞ�	�]���@�؛����,�w�Q�qKaa��X*�R��<:�J�S�`�W�iK���B	�C9�,��������D��'� h�o�TI!/X���M���5z�ڷ�/�Y�qĕ��\�C^�����������ג��$S�ʹ3ل#V��r�O�ؖ�p�w�f�t��}W��S�\�+�7\�N5���f�]�p�"[T�D��ۏ�_��uvv�f������_�.���{�a���W����>�5�"�KZ~���J��\S����^�zspГtGW�� 7;�#xq��7XM� �i��D�F��u+�{��|����[����{��Pp��J�����Z�?��=���4)���a�hz��GD	?ݺP��	-�VO/d*wM@M����
<fBU����eW�IYɺC�1u��S��������5���H�X2y�5V�@޾�+�. l�5�aeƄ[n5aM4�Ɠo���S�q����|�ˉ
�(Ș�����K�Ԉ��� ���/�	�v�+bkF�Q��#?*�Ԟ��vШ�~��|�����xA��R�~�T�^/oQ�0e�����Ƹ��������\�91��A�No��?�bR?]Į��)&&�%���e�U��ѽ��3�2���$�}1�DQ���[��6Å3!	9�o�6�?x�T��G��e`�Y�-+,999_�\G�͕"��.���܁\ȷ�X���\���Jy������Gp��L_;��y88�䎳 n�����*K[��+/S�_���3n�)�K��H�[���?r���u�#���<V�k��s���2�(����B�Vl4U��dqa�3�
f��ʄ�X�$;�',�����yxr�RdY�54�D�>����ׄ����O4ϑ�m�G��"��ɗ���P��}C�Q��sؔ¹
l����A��'ob�pw�>A�q�7��{�8
�hi���8A���=�d���~���$�Y6̄Y���e�^0g��}�-�˸R�ޑ��m	���8g�4�ח�ó�h�3������>7��>�o�9CS��5T�j繐G�B��\�3ԝ�����`�}M�e#�.�vK���*�]�������u8>F������e]ԿC��u�O�L4�.��H�*�nޠE{�F�uӏ�E2W�
/�+X�	R]��K�)�B���W����u�?����7�ӝqoI<��v{�e+�'�x�VU��{�h����=��:�eQWV��R�bg��vѾ�Uh'�n-\�Q�/m�
���&]f*P����8.(�����d��:3��	!��â�;����7X��>r�~Tu�=gb�Z-�>_�["H�n/�a���K�{<`��,:o�;��ci�V`�,�h*�i�XU�g���^�T�bsr(V�D�����U�_p���K��ÂABe����f�:���q�?�V@��RQ�L`na�ix@�Z��ܞ�����g���.Kp����Eb����]+kd�vz�����,�>�;�I����p,��Ç���]k%��$Q}}}���:�5��9�E�������r���Q�t-{䉵d��x0���>x�<K��3v�����0��m�� �����y��䃔��&뢗�'�����i~F9!�UH	4�Cu�1�� g�濖�L��؁��Xy�r�\a�V�Llnn���t��S�N�-l���'hӷ
�� �;���/����!����_�	N
F�zf�����dt�cFA5���^�UfA�Zu�9)i�lA�d���WTo�	z$ ��F��P���n��|�����B`�N����G�Xg�dLyy"�>�wB��߇��\PX�)z���2kH�E��Ӧ�;��#�:���t}�6����5��Kd�����}��X�L`��.��~��P��&=NPY�N�n�,��/�|���S/��g�/ʮ�vyX���]{b�滆��3T�d=<�$�Xr?��CF����gryX�ԙ��i�����*��0��e��\;"�ps;j�jr}Hr��%�6����x�P@����i��=�]��pK[��[J2�R> 0�7�BKl�/��/
�K_��	��t��C�LNNc�c���q��=Q�󆼞��^0��Oy��Vg������ e�^,N�����d����.+j/h�Nq�6�U�&���Z�fbr���`�>�&��lsFe9�X����[����5)����Q#�|h̢+� z=i���3.Z�<11QǔȨ?�4�� me�p�IS��
S���Y ��".`��ԙ��\��ҏv��_l\\���n<;P�Ԕ-�Mt٠S��(�������շ���`N͆�_������q#F%4?�:UFU������rz�]���~��\�[M�n�g���>`�S[[[��;�����Ph�67w��7�39�-���
���CX�3��yh�R��j��H�tvvf�'��X4�<`Jj����H�?�+F����^;pr�����e�I�+<]+ �	�zzzZh�t�B]���@�%SiQY`ٲN�\��R&'ݔ?h����:]�V� mu٢�f�&sh)�fK{�=<��P��-ҐM���N�@�~s�5����qxju�K��h��lv�2L�Y�ͨC���{�3��
9��S ��(�7���_�+oI%�b**-�X��(ⶵ٩I�#\e��d��u�(]PQQ���KNO�+@00�Ծd��|�UN��DGGG��V��.�����)���n�,Z��e�nL|�tG�e��fuH�����8���>`)\�کEq�F�E?�����Ō��f��i��"_���(5��׆<M�u��b�B3���<�C�j}�x���އM,��:r/YF�\"��"E���=�v����|b����R�=�W�ta�޶�璋7z[��~�y�Zٛ=H�^�C�o��)��s���=3]���_w$�;o2p�8������wށ8����GyR;@���v�ꏷ�99�������/�Uȳ��>������y222+3]=��'`���*�����CCC��&�}��:wy�?���9���������_h��K��P6��&ݴ��ٓ��̃��%c{�K"4�Z���4�~	B&���1rUN�h�td�#�GPs�MH�3�%�Lm�jӛcb ��q�t�����c��;��]�WٵJDPWV�+��.J=Ӆ?Z��N�3; �#��!��1N��iN+�TZ@����B�vu�-7������k����p�?�꯯�N��y���V���o�w����bS:7��Im�����M��D�����a�����_OA?*�<;��>�f�_��'?I�x;9�Ư��S�c�Ϝ�{7E����W\��h�	xv��ġ]��rq)Ĥ�9��t�`3G"E��$�����S�!�>�D	�%�B��|]sՇ�<����K���"���k���p1���� ��vK.v~�D���G�OS�ͪ��瑧��9�iԖ�Vw�,,縕Y���r������!o<_	õ<����+��������n�D��7�_#���NC��V��i��|�n�m��˜�6q�&����P���Ē�.�B9�����΋@7�!T}��ƊCW��Z8�۰�&F��b���\���e/�;���0a�6&$�"]\\ ��(,\H�K2Щ=K4��w%����&�%ʆ�25I.�;��U���#=�VB��°�F�^�ТT�"$�z:�5�:$N�8۝�a.��i�n�C�u��!��5���bJdVݥU%R[���s-���}��\6�	��!�����՟�yR��?_5��r'�"W����=�:İ��򻰨�/[��g��ot3�55R|!����4%u����r�����`sV�>�p'�Oۀ��M�ŵ�!"�8w\1`�<�*������g��W#�^(�k*T������}q�%��w*����*ɸ�[�Vi"J����ݔ�aQ��0Y���ɧ�a�E]��Ο���	I7�:�����ܣ�G�(�[_6Z����X�{j��y˗�g�Z�U��cw�:�1�%VI�G4:�p�
�vy���ĕ
+;��0i�_��Z����6�M�ǒ�
/�<��@;�DݶBM�U_ Z��՚Ҳ]�>�2�amu=!;��1�g����/5'�ͅ��"=�s�k���v*���G�c����9�<��?��O��s�d���m-���}zG�e��02R�R��}�*��_��5q4y5aC���G4��R����e���W̌����������#oF0����~��Y��@�~�P�vrPk�V�q����|
ћCB�~Jh��GO�r��-u�PIԅ��K����ِv�Z<�ʚZ��M��8E��v'^�48�@���JXc�	�<2"d+�c�����ҹ�4�$�{W��z���>}hY��R%��5��~�q�h�Q���k.�y5
��wv�W�g����ɗ�%+]"X����.��MW���R��3vp��t��ދ���T1x5Z�h�n]u>D4�צJ�ۇΎ+*T��\9���}���i����|�|����(^���s#Z�5�]�vэ���ĵT�Q��]���-�JL�/u|q��dKn�bΌ=Ito�j�S/k���E�^Ws�:�)������UEBN<��R��z}�å)�҅��i�7�U��o�opq�q��e��=9�NC���mP��o�󸈫0#׮È�O� �y��+�ֱ�/SF9���c}!ޯMרH�`�բ
9g���(�Ό������K�M�|q��w� Vr��$����8i��ܝ�;��W��!���@#~^���
ǖ_2Y�C�7H��d���uk�B��X��,ת��{�l�K�W)k�mPͧl%��bdi����ң�LPDs/GӪ�t�m���m����XH�v]�&����wS��?7, �=�Y�пw�/��W'°K�J>V��>t���O�	Q	��+��oP��l�Ǘʩ.�f^�(_ݒ��͂۴���9�}	��{�*��1ۧ$�g"���XW����Cj���9*T1a�T�]sv(	g��R�¼h��-\�yA~</GfKO\N�y��O�0����%�cɆ0�A���Z�����G|��4 �Q�W���q�������=y��e�zf�I�\L^jG��\B�Y( /�{�J�w,���	o�'���t��g��j�M��MT���m'g*Qs�6>��"�ǈ�xo��:����sTH�W�l$�{P9w�[�U�Mc6�of�Q�𴮾�Qu������_0c��+�/V�����[�9���l��G��5z*nI4ή���l�<?3��5'��:�n���&�B*��e)�	}�#���Zm��WI^i�a��-�+�o��U.仰�u~�;?ZC���Ĥ��l�
�D��#L`{�s�7Ҫ�b�}(�4^k �l�'[�l��\h��$-Qo2��T6��oe�����+����z�������@X��-�8�]�i�\z��`x�3^#�]Oh�u��Ls�r��X����V�#�w���׈�\]e�H8��QMu�c55dlQ�㫧��)�V�p��2k���X_���xZ�o#n�M�Br%�$�ƭj�V�/���r���N��&�^���mw��*/����M�x�c�cx���������7ڙ���.9������a�k�H�å9/�#p�7&ν�c������h�	o��PO��S!�҇Mn1�B�8W�RH���K>�_�Q�=�׍��Z;#���g%�G��l^)V,����-��yiɳ`N���Bn!G}���15/qCy=&���4�����dM������	�{R�f��Mѫ|���u�t �`���OA�9�wh�P��8.�g��{��h͗���Xʩ~(9��*�u`I�r	YTekd�qA�4Ds����ͬ���	�=�nհ���� 7�{���BU��B�����w|�gA�:��D�l#��t��CIw��ê#����β��Ȋ�e��RM���v�q�gc��c4�3s��^��b���h��n\X�@�5&��F�/�5�����S���ޭ��f������=xr��[���w�i�8��61�����!��6�%'_�kظ9	kT���;���plX8F?Y���9��Ԫ���P���)1{��� ^�YSs�B���2>Y�󎭭�y)-P瑘�m�vcU�c��G�x�����<�q���޺T�5I���Q1N������;����k"q�.#�zzzK"���YQtC7�4ٜsaxm�X��Ƌ�J*��|0Io�F+WԻ���z4_b\�����FH��f��������@1��:��j$Y�.��+�!+���c��ѹ7A��!5,AK_]�\�_1�0!�Zc�q
1X[�#�&�sL�^`Z���)kw�E�W&ʀ�WY��h����,����%����j$�ZV��x�$Er1����.���[#ۄ|�(��p�Y%a��Z��DZ�g,`�q�ڧ��.���^t#�m��'\�4�<�e�
4�<ahZr�
ȝzz�]9�)S,c�(F������H�<�-9hX�aA��#��lT���oe:Z ���9)o��f
X��լ��W9y�^=w!����%�O��G-��8L�����ۡ���-�p_�3HC�� �)5v���9�CV�+ҽ[�������2�S�u�QUz=�x^R�Sc�O�	C��u��~@$�ߕ9���<�?�R�1�	4�d����8x>�Cn�xn��l�xt�7�X�#ӷ���Q�Iŷ�ͨ~mw�ʍ;��ӡe� ����_�8C,���$�4(�V'2�8�hiZ�ϔ��� ����]�Xl���[4j�>��]�hğ�,'Ʒ���3E�+X��ي��uu��k%���T�;*�%��#T6A��NC�߰��kZX��\j���NL0��`r���Ṃ��'�@�d�����\�Z��r�v��%o��s6�g=���K�$,�ñ oБ��cG���[�l�<�#x�y\�(��[��j�YR�b������m�@B֭釋0�z�e�j����ܱ������)�f���c-�<l,Fs$b��7����69)�	�ל�3�7�1�T`��]�.{_h>yQG�2���Y��y��.��쒳��#�|/K�]�cā<����y��
y�~�4i(�@bg7�rYG��N�r�զ�e�<��E^�䜈J�=6��E�o&b���C�[_���l�a+��?+��d���v)�r��k� a9=�Q�
t$"��	y���5�g'�ȘU�ѵ���0.����f�eǎ����o'?C1�.j�o�
T�4켒e�� \����3ɍ��4ߚۯ0�����=�Z~�ϣ�J�0���A�E��Z,�F[�P�AU�؁��*;�P[�Tp�����٭C���)��������Kx�\�ĭ��܋\L��9��ҷ��{�Q\�ّ8��;�Y��<��T+�a�ǛҷP����I5`��������A���v��کk/��o_��Ӹ݃�|T�(ˋ�.�'���ߏO�\#�����{���/!�`��{�a=I���KA��r5]"��.�FJƥ����B~���U��Zv�Z»�\�8w ���U���9<h���c��ނ�ԓlmF����	Une�������W�@!�kڂ_h ي�ra���03/��w�����{��U� D��rg9�D�~2x%��������@<��T.�g�%�/L����4�`��S_-��^.T���ު �9b�8��� �����tՙ�z|�A��*r�4u�7g�Z�36�7Ns�]f/KK�X����2i�o �xy�d��0[���Q�����L$Y�JG+i��EP��9t=���r�k,޻�2'�9݋9�W]ϧ�`��F�e�/�:a��z�a��Y��w��5#��6���O��X|6��=���θ
�@��Rt�W6р ��Pէ���٘-f�����bV��Ǐ��ܤ��
�ζȖh��I%��#����*�PY��6����X$%�{��,����R��C��`zV�G�b�:�1X}۞�~5�4)XSs�]~� �|��k6D��,��R�Hҡ΄Zua�@�D��amHUE�9��?��A:�*�hQF����^�a�����@X��_f�z7a�k����ـ����d��D �#�h+��0;+y�tLP��֜��������0���.�w����m�m��}@�>���ʒ�wu�Z1����.�[�W(�l<���?39��R�j�{���Jl�����m��׉�%BCbZ�AM����D��bS�*�u�z�V�q�5MBoRԕ�,{i}ix���İ���~��'┋Ͼ��<���k }�j�Y��WGA7�݋mN��?�M�B���[Z5!�4��^���9���`ԣt3������0�z���a@��P\��bsG�����ʂ�k��H��<٢����`xu���|�Q�R�՞Ae<=3R�&�l�G���}Z�j�M	��d�@�"��Ճ�CE��#��4ݮYH�K�T��zh�[�J����(�p���7R����*��m� ��17M�Z�H�2am�O�����1bq�$mc:G�Ve�sd��."L�G$UWc�5��4��!lY�Ӆx|)� )-�<|��ǝ3"Q���C��[��Lu�B7�6��a5��Nꌊ��J���a�4�3�uQ��bQ�yM�e�����f�95u+�x�����h[Ȝ��㒪��5ԵӶ[�Z'������L� 4)j�w��T�J`������1�2£��uO��Uq�-T���Пcgq�;LR^FA]P�ܝ�Ea���[7��_L̟\hԲ?_m��c��EGPO��)�h/�*?�GF=��6 �ҡ��ߪg�y''?��]6��ز��73���*"�����1+_O�(���^�i逭���/�h-)7�(+�����+;PR�.���Ц�����7m�^~���q�7y�j��X��G��!����?��M��vJ�4���wu4��C�j��2� ��>t��7Q^@Yʻ�ӡi|��v;��>J��u�OQ3��5sV�Z [��j���P(����
br��ۮ_`��vKX�C.�Dc�gC@r$�IK���܊��D i�ޏl��>�@u��"i�/`�k�qg�d2��n�G�j�5�(vv����C,P����Q�@�5��	F�7�k��Ҩ�v�A�?X�vg���/�U� -_Mwܑ�7��op�����@��u��	M�.���<�ܫ���5�)���F�NL	 	�(�F˂�2�q�G�W�4����0F'48���H�`5��V��YTl��[���Tax!Ǥ�)�����R��(���?RQ`�>�q�`�a纼��]��.�՚�p

��J����l�����+��/\�Ҿ����L��Wy��H��Z�R�������J��ƨ������v�+�[8U�V�Q��)/!=�5ש��N��;ŧ���zm.�L�oB�Ӊ+�f�����A�l�,��3�i��ã#��WR�>I�3 ���9�$�h͈��O��j��VZhC����^~U���U����ZH�R�3曄'V:�iW��}&�Y��Y�^,�,��ʓw��
l�L����G,�l�	�1bN��&X���kX.�?$x�@b�%P%]�TO1�����P�ˢM�k!���[�^|�;<�I�h�>p��͛�;�U�RKv6�ޗMO��yj���%�K�.cP��k���
���X��]u@P%���c��`�P�%^ JH_�N/�f%�i�q��Q��,O�q������+Xь7�/}��3A���iɕGF�}F����S��u��rer�$y05E���kt�'MF0���l�F�N�v�p5�l���.0��:֬�S�霐�ˍbz[��bH�E|�^	�c]�,P�3����6:��R�ԟ&=��ZF�5UC<�֯_��6�Ar>}u�-��1Jڇ|�㿖�k�Ԣ��ÏT[}��&����4�&��yR�;}ݨ��*�Z[�e�!<i�+P�P��^*Zhw�.����[�f�M�識�1A��r���O���T�r8Y}�ՏP
k`�@.��q��z�U��(f�'�/y��<�_���N E @i����J�אռ����K��H0�m��x�����5#t6�L�
V�淐����8Uc
�8/�	X�.1��h�%4�Eh���v=����g��2�6�Թ�q��=L��j�FOC��4��N�Gծ@I@�@`@]ZI�@g�ݾ�.�R�F!շ��V�=!�#@�^tC�����ٍM:����By��$�O��(4h�n�"F�M��N�M���lm�[E��z�:��%��}Y/��ش���9���R�H���gh�!�t�w��8�D�fc�w�q�hrv}���8�Tt�q��>��V�S�>S+�k�	�Mvx�7֥`�Ɉቘ������Q��U(�!�I6[��]��c5��_�ʷj��j��+-�ǫ��9�.>�幒��s�0�YB�JU/�K<�ڄ^{{����(���Z���4����P�M��\�`6�OU�R#�.�+����©�c�%WS����,K	�m�C���L��U+*	4�O�Z?�|�8��_w�
��+��\aD�I	A��������ܒ��|u�E~?-�Z�Bu�6�A\������H �/#s �W�ďjjO�x�vO��k��7���4�	���C��ayD�6���Y�d�����'Y9���q'p��z��B�i~���S�g�33�x�T��%���{'�!j� �O
��9�4�l�B���Q��V�w0�`���Y��eM��٨g����Қ�Q��'������^g����Åѣj��K�=��j�#HS�����"�!�+�;�N�`W�U���Ĉ��D'���-�r	@�ԓD��gG�B�\yWԳ�t\����s��~cE���'*3!ސ��4�pѤG1�8u�^���P���!��e�e�k�a�9���þ��l�~.Б��zFZ��T]i��+��τ�|�
�R�I2alY�_�'��?$1 dI�92n|VVǨ��-W�L�p�TT�)<��xT���]�bƆ.�B�JHN)We���{�%򬩥�i>^П�E�a_�Ɖ,�Bi`%��ƨ��U^}S���oT_�{��7�J���-Z3��{}�CYAt~!|��Ja��`y�`�R`�S��]3s�$�(��֯_>�6
!Tױ5aa��1�4ػ'g� �t�_̛�=�����v�u����v����gl@����1��*����ꗆ�M��0�[-�lxA;\���`ݼ����1�|p:H�]5��y���yŚ`��GkLô�a���O��m�k����13JқC�Z0G��RG��e��������D%Y� �77���gxAmWk�!���/����g�s�b��8W�|FY��7�%b���
����X%u��>,�֍�_&:�7R$��zt񵒊
g|�u�=䒾/=G���������Wm	��=�ԾR���RB/%;�d$�r��s��JO,���澄��ڥ������;F�`v�������/t�j��+�a����{���_\������_�����g������V�Ż�7PK   6��X� ��! �3 /   images/199a26a2-2ca8-4fec-b52d-fcf4e34cacf1.pngd{eP\A��������݃���u��%�BBܝ �%�Kp�`����߭�����vg��������5�1���@ ����.��!��B�	���TwC/(���.��^�%�����7[o?O����������������	2��� ���a�A1��T=o!�Ŗٖ���A���GT噧cԅr�k��,����vH58Q�ͤq�������Å3x�HI^c�P�~Q{��gxei{�v�Jv�"�����pI��í�m��͔	��8�g� ��v)�Ep+uc�aʪ�b	D���� O��8x��A������#�֟���OQ<#�����F�[�<Q�kU_,j	����},��php��E�l�z���:^)�����z�o�FR"��:���y���B�	��.���'�җ9����l�휗9d	>��z�w�/s��#�Ү?��@��C�]��s9�����D�z>�RF!�Xj��h�G��rѩg[xq�h��2�i�����$id&�`EQ��R,楚�Pĩ�W^ }��ƽ܅c��??���`.q���d���/*�
�9S���L�(���{���8��j��ѹ���b��Mҥ�����U��#I���ջlA���G�,��ϐH)l��̑�������Ļ����Ĳ!��jV�H��`bG�ϻ�2.q�",̮����H���r��1#��OVp5�-A�[��%��q���H��]���<9�6��&EB�(R���n"0��_�մ�9Z	b�@���&�ghk����������.n��x�}Z�V����!���UT8���<<
]�`����s�ǔ���{��x:_�7�K�!���B��Q:9ځ�)��+Gг����蒖t��d�E+�^4j-���?�|b઺=hzQ�w��)!�nա�9��
�-�W�_kVg��Qe��7et�R����edע�g���T��{T�q�O/dՐ>�o����5c�,�����}xW�$x�)o��_���ƈ�8�2�z�#��7~hP��4�h��}�/���'z������و��ޟ^r���}pCY�E��~� �p�J���Q��[�y�f��� q�+FO)#�$���9)�Y�����������o�*�*�����]�{�3���Ji�<�e�y:ɣ{��U4�bf��߮	͛ͮ��e�i�<�#����~g��Ro(�8�EA�{�`��A�������ټ6JńY�-+��+��ȤX��o֚˙���6�J��}�	�`B>B:�_uI*	�����VB_@�q��������r�����l�����7�t�<�D�ë�uD�Hw��jjǢCS����t�H[`}KL�O�38����݇���R@AzE�h�"��n�T��Iy�.���.���^y
?ܲ��f�;�i�3SU�N�Ä��	��{J��� �z�@�������[s}{]�,�i+E`ЙV�:�y����ïH��wy{)N�o;���^<l�~Ic�
�������w�Z=%�^�X	�ů���NWD
�j�d<�N-ۮl�
{E��������|����=���?}�"�$� ��#���(�vG"����
��P��?D�zr ��j���`�����l��0e�z}�~X��q��S�i�Qʸ���A��a%�;>�l�5EG`���ul$��̍#�EOC5�G�>}�Br�0��8�"=L�o�]x'�^���wxz��~�S���.��NA�d���Z�p�~4��Y-Ƕ��=�L��q�̸WO�s�*{���Qf�)%��H�¤��:���� �K25��eË�%y��@q���	K�"�ŗ�c�/���4���oxY�[�	ت���"}?>�eF2��(*8�@&	|���%/��b��$�m�
@V"�83�`Q�������c��D��Fx^,g�WeN�R^M6Ŷl �j&O�DE�^���� ʍ�G����s��Ʋq��r��xVa�*x=�^�pEt}��҂���k�$/�� �K+��v?I��$iߞU�M���2�;�;q�1��b$��a�,��[څ�f[c�Q��Ř�(�c�����ڲw!&/c�3�������Tm�㉗����nW��7����-��r瓚'!�`B���
���>Pb�a!�������M���p���u/pz��Ӵ�s�'L&2�&�R�MY?� ���B�֞>/̂+�]�����`�R<va�LZȟi�*i=���)z����ē1|Y�D�"�QA =�3�`�2�b-�����r�/Y-	G��tk+h����^&Z�b3�I��/�M�@}uf/�ሺ��:�b�Y��x����ǳ��զۭ�^`��<II�L<�ۖ@��z>wD�:I$1((��{������}7�.6鯿��XdYX��J�;���h����0�1LO�78
�����������5u	T-���?�œ���Z����Ya:r%��<��W�S���i��e�0�s9�hi��I�)���OU��t�u���6x���zA���}��l����d	�1��ˀ��7��^����S?�ʺk��O�bG�����3{����⬰�pQ��Z��'�7�s����J���=������m����$�Nrca��Bn����٦4�cЅ�(�nTTACz�� bg�ϠU)�n�2�g�kƹ$��_�ߠM͞��T�u��R}>!�s�U:��9�����y�QQtLEc�wT+,����W��s�7��4v%:#JmiD�ٕr�2��S˲$�U���E����5�C�e+2���B�&��P�?8q�ʘk�`�0m&9����9Ë�Zﬀe'P{Џ>�N~y�aܑ�,���h�>��cY��E-�D�x�'�Нv�O	�T�u-Q ��$�(Q�4-ZI��ړKI�J�ײ��Jr���.j�Z�L�#~%�J�s��&fEyq��yjB��?rO}�i2��������Fz��_o��(ŠId2;�P����q��@�Z2&�ؓj�F�^	s-��u���^ �xG.?��d�5���W��+�|��-�^�%{92'��z���K]V��O{ou1�N� *�,
�0~Ca�(%�?��-fx��*�b�= ��i�<M��Kc�z�J��b�'���Mw�d�3�*@�&G�_��*jW\�:�W�z�"��hF&�--�^�6:p�S������ͫ�N։��KL����L���e�R���2�� �GǸKǵ�^�^ u�H���EJ�#�����V*�	�g�m�����9���"\-���%��d�/���#�F#ˋ[6����t秫�wf�ӮTF�ߟ���+�G����H�`�mW�9�X+:�K�25풮���_���8�a�
&�G0�Ac��.hP5�_X�Y���b��]��0�޳	�K�#a�54K'�
 ǂj-F�}�z�
�totIo�/y����b��5��!�h��T��D�������N�݌�r����ԛYOʸRnIJ�ym�-���g�:�n�I��.WU6E���;m������6����T=Wb1igG�ԍ�~�h�8���}�����D+	�#���Z3	�w͒��U�^Hc ?�jn��p ��|#������% d7$�Ю*ǝ��4\)V?TP��PbW�mN<���'ؑH�ZbջH��,�i�����!�����]���� �c�3*��Z���tG���pؐ33dS��Tу���1��s~�>fd���+�	����_�ӓc��?�.���b��УA��;+�����I���J<��am'La�l��������;���dͶ�!u���
x�]��=sSq�UVi�Qb_�M3��Fv��t�6�J�Fv-���fki�B�('�Y�FJà��s�kiW���P[�p?4		�Y9��.������֙x>>V1�0`���TNLSd��y�0����!��#�v0��E��%<TK��,C��z$�6�}�����V��A
W���y��P���������W�G�2'r������Я!�Xǎb���o�Wﻈ��1FZWi�\�Q��_Κ��JFQ�{�׻�:Q�܋�>�?ny�"*�U��#��?��r�FJ7Q�D6z��5���()��E*��708�J�}?	�`:�O�4�4}��1�� �F����]�@�Lͣ�L��ۊh�����|��F�4��ݥ�����O-����-��誰��!��vOr;͇���1�0�o� -:�l��\d!���+'֗O)���wͰ$�L�S��Z�,��/`���@��{�@@bA���9]��q� ����Bˁ�7UeݭQ�YG���s��=�J������GN�w.�E%/���v��/����hʡ[�"Ek՞����Nt�`�
D�������H!�GO����S�	;�UP��t8b� cL�A�=MG���' ��T��-KH��KG���:)e3Y����������Xw��mĆ�����x~�����<���l����M�}��\�`�i+��M�gzu�]�ՀA<��Ԣ���O��4L��⏢����cɋ��7�$_%���W�
��n~Jh�/:H����|�')7?���'@�|JR侄)L;����R隭�����0�/��n���W�E�ܢ��&�E���{�Oo��|d��MM��'����\���c�H�#�c���?<�2�Ua(���}^��"����>֫�����U�k�nK��l&�K�ۏ�F�2�fc��$Ǿi@}�c܇��.��)��I᥃��И�a�s�-������ƿ0���9��ó��_7e �rſ���!����U� Ds0E��X)e��i���-�8�b��O�؅~�1"Be%ݼlD�\^��|�4��E#���є��uV��"f�_da>���3�!�8������|D��_;l�"Ҟ|�>{z��m����I���i#�(Mx=�5��рA�Dq��?����7�y~.��C�����!�j�q=]O~��^�}��-�L��eaI ��.����{��sH}aB~"�r(t��=fW��u}�z�{f����t�΀F��r�ZHWtB>s�i��#�b~�L,z3ܶ�|31Y'�x�k�:m͕Niɩ��)�f������O�3��o���I�"T[�J$���~U�oh�B\�Vx���X�����LK�����T���'���V�o]���܂�ECM0-zS�d��EM��c��â��n�U�A���]�J�w�sg�C�}��P$l��:�n������U^Z��P���&���o�-��w�6���W�Y�Z����|�jU<W�|r��:,�B8!vcբ�v�#�		�d�a���)pۢ��񟔡�_1B�&~���e�shF��.�®+��!|B�y������R����/4�L~Ws�fЅY=��3x�/��t������߇@_��kv���{�����@X�˟|���H��1����
w��#��ݼ1f���Đ�dv|i��47%x�������A���a�=�K�E��\���Y�?�m»��A��ju��Y�eD�vE�~���&�1�ްXڏ{�s�tD�y�ῗu�mK-z��廪��ɛ���L���2�fd���Zb=3^J�!����Lzc����#���	C@�B:��η�Z#q6�T\Z����M�f�Z��υ��nd#YX�$�󀾣��V1Moa�<PB.o��^����%T^�ڣ�JVSmC��P4�*��󒿌�^9A��Jbw^�6�滚����]��M������4��A��S�y�)��.�����j�+֌�2M��*L���X��_K�|&;�^V<��,�~cͻ^�}�߇����53��P�ճ�Ɩ�E;�8����Sr�KJX�\����.-g����i�4��Tp�"��@�M��)K��mR��(���I�>��]ރ7��?z�>8T��a�N}~���HU�Jh�WX�a��LV�C�-Q+&w���x\����[��b���=|nu[IFӒ�����g�q|/�n��G�^�	X<|�b��o�w��n�'��8llC�h�����I�� #�Q���`�����Ev�y�̫�=��v~uRBu�-\z�$�zf'!�ی�KP?rZ�J�앯�w���k����yH��'��K��Eќ�G�H����@'��#&�����'�R�.��Lb��(1���)79�aq�!d���`!�m��<��S�ו5�dO-�E��\��P��4:��O~e��^�͏�Z����x�pW�]��p���B	������-�%V�*�z���w�����iiy��{�Q�'�c'*���W`2F~�w�]s��`��? ��8��+���#����~GԷ�L����fm�ݝ�e���C�[��4�_�����0/�Fxu�<j�������Tw�Rf^��i`4f$ ʎ)��px�CNW�)�'����"6� Y�� �P~�,�,����Ik|���I�0]�5 ��҈��t�d�d��m���<�q���C9�k&���;v��K
�Di��	o��Ĕ�;"t�̥��߆��`D6�GB�R��g#?���0-���%M���c����8N�+I���FH�8��M���QGr��1�9���M&4�|��<1\Ƴ��S?};�(T�QRմ��������Kj�<UT��w.9��Ƃ��W]|s���մ�`�ѣ�ܨ��IB�}o9��}+wa ���)A&e"��S�f]^}ɸ�'�i����kw��4��Sek�L\�_1W6t�Bo��_E�X���~'����=���>d��$�C����т��uj?�KOԬw��Q=�I�H�)����4��k�Snc?����0W:)D�Us����.���T���L�Ј��א_�`�x�9U��*��?ކ�n'xe.�H��IbG�bV�Y��bw%2�`ǝ1�F�ڷ�����QKV�
{xd���ț���Z�<���\5�����oY�\RWry���J�UT �5���X�EE�	�ӫ ��C��d�� v�?�k�%T�bu�����ܪ�� ��*E�4��ߑ�]�dIPۥ_N��X�񸓼�n8��6��7�K�j[�G�B�]T�W��N:�}�[�*�1�;����Y3�;��.�Ru뀟�"��~-3:�ug<��g�L�#�I������r�C��"�<�z'��뙼�ET�(g�hP;\�8�q�͵��9 �%!�Y�O�����W�I�0+�"C�v���]�K[KLܽY�h	ie� ejf�He��������[�C��]E�� �99�>#ۍ\���tq��fW�#�������p;�[?蟓XmA;F����awjM��w�A���+t��!���Y���nץnt�!�1�b7U��c��.��<պy6�)��3�giQ
���T���+��k���J�v� ��[���Iǌ���!�N{���zQV��%L��^������@�t����|1��� ~a�}u�)��1nt=��2�#��N���6�9������Q�IDK��\��������Pǭt�η��}��v$�_�[^v�bFKk�Ƹ($���ͧ��e�'�6�x_��9�F�ږ���,/IBI;�lQB�N>@�U�ȟn�i	il�mOL���#u.��[�^����:��$!���^�q�䭭Er@U�P�+fʡ�/��Ao5Y���	2�����p�Y8
c�#ؼ}�h֙�bH&�p��ޢ-���O-Ufs�G���-{�8�M���c}"T�d���} 6V���M��u��H���Y�=13~�����*�Qyu�v.���Կˋ���T����D�����C�ώ��ꂴR���>���c��]7/�e��9��L�g�
Z��1�h$�q���V}1�60f���I�ۃ�=37}����E�vtT�W��Lj[�HY6��f�cG��f��=x$H�La��ub����.���y�FLR�|�N-=��v��_T~?q'��9GnJT�޲}��D$��m�rb������v3149�(w��ܩiyV������Y��P���)��RĮ��*V��[��_7i���8E揷�ڦ��$���(�@{l�"Z�]�#_'9�lO�o�cж�T������gs�)�LH<ұ�����g�����"X�,��Z���E������|��ղK��0�}	�17^�z���mVq�!��?]��W��2�rhT��Ր#�`W6��TX�Ҧ��mZ��ƅ���cn��Վ�<��O���r�|-��,[�,
6Hˠ
�#�|HN�w��W����(>�-H��{��c�%L~(�+��J+��r��96+(�	���hל6ͪp�H�{��{�8��E��B\_(����t�*{n�6�ݫ���
91˵7�Z���E�6����ܦ�?g��՞��j���PY]�~��_@��囬���̒�<M�{D5��{����J���[� �!��7��񛔏�c�ba��}N�)�����j�G鶬�1S�٬L�a�%Ҙ�Ť����\)@����4��������lV؍��m� �E�"9/�K��b�eC��K�qw�t��}$�W����g��{�����;����x_��'kf}�u��e����1�U�篆�k�7�|<�+j</�I)����P>d\�����	����ڧ4Eq�xvW���l�t(�z�:�H��=j����Nf̉��F�F��͇��o�!C��q�" �'�����4�5�[S����w+)�=o�ܔZ;
�9�Y�Q���G3����W��a�PV�	�@%�z- ����&¾�gb���*g�i�'���$#�i����_�J�|�u�;��r;�T��G�q�u!p[���v0���ܴo�%5�8P�L! f�k��z)|���o4c��c?YP
^����M�EHg7�o�07y_���2Ƕ��Lj�w�S��m�0�_�Xk��DǴ+��v�
���m�KO�<S����U�_�o�3i�FP2eO"\絴Ay���0���4�86y��QW3	���J�s�zY�����8*TX�������0=MG����(��(#R�q����a,���(��۞�}�0��6�wC�ߖ��0�F[���(��ٹ����b�'���j�[�y��k>���Q5��mqVE)��:!sC�[�3ʸ�_�4u��K������(�C���`j�V�
�����J�4�������<~�O뾋�cl�v�Xt�N���~Rn?���`�
�RjHV%Mu�+"�2�����d�K�r�eF�)A����nL�5d6��q���m��ʿ`:����N�g@Q�nqF��J��}2,�-p���F�.�t����^�@B�����A3(�������j�6���@��v��#�Ƚ1�T��P�J�q�a�	Rh@�k!��mNR��*�V���Ns#�;5T�K��Fd����b`>]٨(��5��T�*����;���Դ��.�V������:����#����vO�1C�M͗���1�%R_�O"q��;(G�J�5���c�y�1
"�ԑ�K3���]"�F��1��gM�f����E����[^[������xݾ�z]4�n��������enNB�>'!���KԢ3��n�5v��#~�L��aJ��������R���5�[�^��Ư#yJ%փ��[���=[9
��;�i&���赏(��>p��,�]vV(����DV�kC_w]&�!��.p�8��8`��-Q��vũA<⢨Ǻ����o�m����=�?�~f��2o�+Ĳ5�ب>��`*K��~��X���m;�ʷ��n��Ն�6w̩���a���&e(�~��s���KWf��0��ϧ�RK&�2�i!�zڊ�ay�H���\�R5k�Tc���Ц^	",�,�h<�0�7�����}�~/���Z��H&)��5�IY�
��� �hDY�F�E� ��;�m��`1��⌳%�i���o4}x~�Ti�2.�)D/�]�U"��(8 -�}�\5v���i������:�80�,Z����	�+oXJ�Rs'$�;$?BE�i��y\�ZL���ۿ�������sn%9>�^����p���kt�����M��'�₳���T:�~R�Jz`'$ŏ/����S�	�9���=�{*a��+Sd2���S�Bbmc�q�	�/���*����k�x5��%_V�>Ӱ/-�n��#�ɠ�R�W�6�����23�9�l���N�e}x���E�˱\�,��K]����YG!Ʀ��آ
S�xu�H�-Ȫ*�!7�L�����^��
��xS���PEl�Di�
�L$v�N@���592���$%EKEIדi nxC�pϯG�~U0�)�"�me뫪���T�2=F^|������Pl�������)$�^�!68XL���!]���N}\�j����"���0qb��T��K";�?�����E��Q�l��DĲ'�pމ���v�*zH�n�R8k���n.e����%3O�(��]�K$�8���`���@��X�嘯���=v(�44��3�<�q6��?���]�:�M�����#�(�_q��0"�p\����+Q׷h)�"�
Jf�Dr�B���J�Q����x]2U�zUO5��s�
���v�̣6��m��5%>�BA�m�ه0�*�pe��e4-Ҥ���RW�U?�DN�F*:U$󎜠��(�?aj/rG��dۊ���)�Ψ,w'D��;��Kga�i_/K'Vx�A̪R�����9��J8���Cj�]�^����|q|�����N��5�}�&@/�M�"M�>Y���]�Z�
�V�ZU�A��u䔖w$�$sS虳'�/C@�s-�ȣ0p�Ԋ�H�6�q��ǩI 6���QW���"�	r;�}�9�ϰ����(V[�YG�RZ�K|���%~?Ib����@�*M���㊭�3�iz�]"��:V�q\J�����al�t:|>�8��V��A�u��<�$�q����@ۺ�
��9����ީڈ֐��OQ�~&����?!Kۛ�0zg�)�n����`�Oa��
��n�O��}��B�?6c��G�8���1�}@������!�9E�e����|�4
$ݲY��j�D��I��@��K:ڱ��0�5?F�}|�����#�k�a �p��x�;d�z�<Qf�O;J�| Qj�
n�=�kOj��.���[8Yr���(��3��&L��Я�_�_t���T��L>�rR��'���ӫ�몢�4`>Ja/�GuI�A����B�S��!
��!2wK��%�,!q�ag�)e.������׆@�}չ�T�nY�a����7��oUVGl�ӱr>^�T:���O��8=/� �78�{׏P���:�^i�K��u�`޼�*[�*�����t6x��d��\�WQ��0��x4TB�C�P��[*�Ph0�_���o�g�@4NE��*�:!��6�=pVLp;�����i#9�!RB���!�a�lx�g��Hf���J¹�8����L�e�ƨ���i�D�$��gQ��r� b/\�8b�-��)�.�!Yޑb�~�Do����3��?�Qhّ� �' �a�t$l-���-��HB�R��T��*'�p,�^�]��Θt:��-B�rroMd���s�rãx'�~F���`�S�"��͠���)#L�?%�!��E�E��Y@�)�<��m�-:���>E�z���̩�N#���A�ސ\X�-�KBTga#$���V�����f3���Sd64}�v�k
�29�QSҢi��e�:z��B惛���ՔOi��

Csl��9XI\-��̧N���e��1�-�oZ����A�Td���7�+��0zYn�/c���&�48g%M�X����jԄ���=ƱR��d���ypS��zHd���+r��Ƒ�̏��|fƍ}�du�~}c���&q�sZO���G���7
���S#t'�:�ہ<ǡ���-�f����8�!�	x�\H�<��0U$Y[���8�k&��z����գnY��R��n�f�Kjv��wh����b���֏����(��/0[PB�)���%>��i|j��BJ�k�sM͹���v����Nj�s�/��68�b��*ѱ�!L���Bt�}iZ��n���J�W����v�|��㏁���K�"E�M�LT�5**��������]����;<yVC�!�����7�;�@&'�v��s �U�7���9�EI'Vj
+!HUYZ_�$���/��:��`���[�~�MU��U��K���f�e��vO�!S��/�N��6܋s2���X�z�:���͚��3e�':�2)��My�y�<31�� x�N��g>�5�5�v&��_c���0n����4���4?i��L�L@��\���	`O+̙��H����B� !��m2ݱ߈Ǧx]��X�Ô��QA8Xd�d��g��w#���޾(Z�IP'��ܕ�Y��՞cv
�A�yq\���
� �wb��=�L�I��y� ֩��e�� ����
A�3r���"��S��j���
�����W�9%B���^Y�鵏�Sq�HHO�����Zx�Z��C��I���D �͈E_l�S=�=Sx�>cp��|�h�®�D[�=9!K8]Y�F�� I�-M����\u��8�h�wЯ��B�|���ɭ���D�ˉ@ 
�3f�����1(mO@�ĥ�����ئ��@q0����E`1���T���L��qK��`\��/}���^n�` ���i��8BO�9��Ht���m��%^�^ݍ���j,"�	�+�C1�� ��~4���J����D��Rrʋ�{XM8(�f��|W��X<�ߎ�N�J>��R^"d�rn�n��;3��(ʞ�Cy�K2�Z7�I ���#�c�L�g`��#�kݽ}�`o����#�G\)Ξ���"�������'� �j�G���S�_P�#����.q<Z���џ�Z���dȰ9�	��n.�k��w�%�sYn�~�-Xrs��j�M����e��A&�Q��1f�M?�=�J�� p)��9���IV(�b�J/?�mŮ�J�6�iҒY�g^��	�/:z�;{g�74���æ�q��ӼtY��4��hϭaI�1��řD;w����?��a,۷�V�,�ݞ:�;�q4�T/}�X���Q�+`?�QgdoJ ����_�Y��>/স�Ce��iդ�����0��n΍i���ز��m�*�UQ����q('[����|Ӄ�f��L>��]�J,��3I���S��fN4�Q�<M�A��[���V�����L^|��� M~-˩b�6�`�ɾk��R
9VE����a�9�,s:���H29ֶvP���0>���ۮ+�s���;�ͳ��]�Ԋx6�<_Ƥf�
���-��eu֊%������?�A\j۷_��K���D2��W��.�5a��%EII�]���	�u��l����xO�{�|�KM���ۤ��A�>V����h؄Գ��Q�r��uq���`�n����]�g���_G����������<5��ޑ3	�(��o��G���(�uS9� �����v���iY.f�C�Z��z��h�=��4�/!|$Y|�\1�l_�+!��I�lp���]j� U,���E<z��y�P���}c_��Xo��"��R��"Ķ~���,}�J�ː�k�nl��f	7����-E6mN)P������$ F�(L*v�T���w���0g�[/��U�E��h\�y؟R�Ս*w�T��������};+zF��<���JBMޛ|S;5���f򥟈CFnCH�)8؋	\��&X8k� Bk���l�ec5�{�r���{Qek�hf��-!҃t %1,9/�ڈ�{}�6T�!I���JxY�C�����>�����ֱ�sts�遌
�H�c�5���I6�c���G*t�lRՀ����q1�d��*�:���ⱈwG�2�ȯ��D&��Bs��Ӷ� @��E�����\�?�F��w���qNN�R��>��F5ل��<�|8�Ve�fHK�1�:Ǵ�X��"j��y�����B�k��&���_�(�xAE�,��NC�䞫02��|w3�;�Zg"�Ժ��kQ� 8���xA���J��=�O���Ob�zst�2���4<�ӧ�v�VH��3E듫¸���&����=���[S���f��an�-��We"|0�6S��'k��oJ!}E�I�$3w/�Ŵ���t�a�;U�?��Y/c"���4�N��op[��~^�s[�����n�8D�)�mNߍ)�9:X��Y�Q0kC9[MT��f�*���;�joUTQ����W�X���8p��'0�$˫%�d	R_��<��6��c��\)�l�I3gn�(tf��!
��j�jI��(�~��4���]����S�)�"WZak�a�|�����Uv���'������c�(�CKNP�/�[�;��ə�5�@i�Y��'�F�{]�7Y���l��������\I����!�N�L(��̥l!ϫZ�W���;�@K#L����7]k\�2Q��$�y��sZ �ȅ��Ϲೃ�Kk������ҊSk���c*qa�U�j9n��ϖ��=P�u��b~5�[�@+X��|�|ۡm� qx�r�e;�<��������o	�+�:1Ӽ�ӝ��MS`]ڹ|�u��FB��+��)���7�C)�����q�K͵17?��X�I����[����䭣���]L��k+��M�'Hf��"���Yq���Y��/�6q.�����E�*;K�LJ���߸�x�o��u[8���<X�*{��H��J�.����=wq�7Ҫm���h�Q�(`���k�@n��i{5�n\����[�Kfa7lg� �MVU�L�ʺP#ޫ~xz����e:�����)��w�f�Xd�{�֍C�߆6��i9�-I�te�fl��� ���0��G1����A�L��H~�0�V7��޽a��G�s�Z?��Js�	�i:0�&\�{�~s�i���d'���ī�m���?�2�8���K����O,B����q�)K�|�Dv����Vsd�w�"���]�u�26u$iO�,�y*p����n�݈�b/���p�ݛ��µҎ5�Q�d��V4��D���b;�9�E��痤נM|]9@:V�E>��S,>�x�	��&]���C��8�dǑ���|P��`+?@�1��S�Ԑ���`۳�6��/�����wQ�5B�p�-T�q�;â��d����yս؂Ui$�)V(1A}4=����.�,{���t�ƭ����%�Н��g	~�L��	��+�^�9�ןo.p1��@C�*�b$��ς��B;�ՙt��7�G�G�ϭb���/����3����z���@�&��\���"��"/`*Q��Dy�]�艐�·�M-u.c1���ԁY���v��P��0��	�ID�j��SD���	��zy����
JY�!�v�#$��֝;�5�Gb�~V�{�����,�{w�s�].��>M}�e|]I�h�\���i��9{ ����-���!S�g����'}Er@�^��*6௯)� �vO�/��S��S����d,s�bt �&yc�hH&$�h�,��t�=���R�y{���f%�m�fh����=k�z�wH�W�F�@�w�,����/J]0�۩��GP���*,R�Ϗ�G��I�����9�`,��Ѓ��E��Ϥĳy�gn�؏���+³{��T��޹#b?�� K1Ж��.!����|7Ϙ598�[r9�yU�꺁�џ�54�L���݇u�I۱�<	n�6DR$5X=.�>��� �4�Au��懎|��V�+.�s��6t�D��,�p�@��C2�bj�C@��(����`����y Y1���eim_g&&0��w*V鞐�?���_Y��QsZ6��|�T��u��_3�_�K]x�G$�g6�8g��몎ݯ�#�J|�.̯�Ԕ�&������X��cn�'[�G��J�N���J[6���_�$Lo�>1�J�;���[�/�$��ZL5��
�O�,��RP�+�s��y���y���9z�lVr�G)O�T;�B��%BOM"O�n���N6V㈮��d��&�k[b`d�����ǳ�v��B��Y[��5՟Ȑ�ˉR�2�E��U}d��	�8@	i����2��B�N[I���=a���$���S���.�W_������b��jֈsb�]_]����f�s�Ur�dr=����³S�k`D�\~B���Y	����Hǜ	ъ���aL�s���#-褕�k��%H�Խ&%��I���#�K�
U;t��Ŝu��*5�<N��r+D$C=�������y���z?�#dP)Μq�K���J�8��n��ə�N�4�������5�5Ì䉏 8ž���n�o���ܕ�	6R���� ����~|	��C)š:~�����5��Uۭ&QqZ}���8#k�;0�H��������C*�ﲾ�CfQ�vkC����"�gY�����[�E���CI�� "  �4�"��"��(% !�]R���H�8�H=�5���;�}�s}����y��b��^�Y�z���g��'���0��f���:w�tg$�	fV��?8�q^p�/^�f�ym�!����/K�h����-�*���^]�l�q>�Rܲ�����a�I�¡|dKT����������)GQ�'Z�X�
�aY5��Y���QV(}˝�{�5)#�	���k����E������O΅ì,V��F���	[^<�[=͒a��ǜ�x}�O>��̞���}�y+���_i���� xI�8�Of^�=��R�#����ƛ��G�9dD�7`��z�4��8�3P�!�Nxވ��/R�>S����+$�� �.ġo?<�W%	ݘ؝�~|�q~*f������p�Ʊ�Js�M�s�4��W��\�+7B��xc��婙���3J1�����=ϩ<��͍��,�!
M)�'-���}���zu�9�?*�q�x_��D�.�R�A.-7�$��F�]�CU�� ��j�&B�C�ӓ@0J7P�=�+y�M�����I�گ��>5������sx���������;տ\-�"@�k]&�^���!W��Aa]��F*�]O��T�����:�����ٓ�����k��4�}�
�r�r�zT�G��/�d�����WO�i���~��|�<�v�l�?�-����w+�i�]�=^�Y�Ԕ؂`��_��_�<�<���Kq�����>�dm���h�C!�u��/6���gM�Y������`��������}�*G�.�|��~&��u?�MG�R�����J��#x�z��+kF���k(E��<o���_�:��x�智�e��ҋ�����������i�N��g��.�p4|����g�C8y��m��k\��oK���wAB�<�Ql���׻h�3
�����f�3I\�����DLǌc&���:�>7i����	�O>�i��9q�A��Z��m�j��ǴRѶ�$M�>��7�'\�V�4sW�-��!.Fx�.B3g/���~��d��[��!���9�cZE��:RC��8�o?~ӽ�����s��g8��C�[�2�4V'����u�i��.�\)��L7;±!3J�>�jU&��^��=$i��Lw5�_��;����qr��s#u��]�m���"��U����^�_�mb.P����������+Gh�;�%�L���Iy�^Ȉ�v�<�Bh����~����諴\�y���܇��a(*nrc"i+���2N����mځ�	��;���q��^�i5G	ߖ����i�A0����1�������;�>�^^<���G��x�
6kZn6����E�}^����H�P�>r�@f�
;D�gԕ�9�>�dL��#Q�xN���h���W�%e2[�'�>,�g,��
J;�ӘG��?}r�N��0�AR@�Pa"����)�)���/�*ve�P���2w]�>ؙ���]4�M�}y��?�e�W��{���$�9^�8+P58Ny�>��8�j�t������s��JR��I[�����E�w�^��DA�`�v��p��Nwb2��P�����?I��=�ťxwf�}����eTA^�T�7������q���33����x�Y2�� +��-V�aՇ$_p~*5�e���uw4p~~�_v� 3d��B�pPk�%�\��T�<����yL�0�J���]�L,��zDH�ʚN�`�'�G�Jc���IF��3���x2�+�l�`#�~P����U�E�'_OeT��O��A��ʬ@1����A~�'�I�f
!�n!Wt:w�c�|7��3�!�+
�z(sRH��sS�>~Od����x��d�����su����\�/��f,)�ψŉ�H�*��o�u2l����������Ē����u�x�9xe^_Z�W<#�S>�{�G�7`�_f3��ə1�+_��b�]�7������~��L����`�9��[x��Fő`���ٸ�I"W�p!�gx�Q��=�Bd�~�퍻����|�t�,��G��fV:+��*}�U�=?�!�<�	l՛����BaQ���H�Wrи�bd�<e��ٰ�>d�Pr�q���}JdΣ�w���D��C�q������z�~������.?�x�<U��[�W3|6W�RCX>+8�I�ֳ���b��Bw�^�$�Ѯ�t���7yQ����������*��1�5x72
����v��w��;SN3����}R�*]�Е�ӳ���+z2g����E������׫(�`�kg���+�"���0u��%ٺ�u[Qˡ��ʳ0*���j���_�A��'�|_�~�1x�Z����R���U��|`��>u�Z8J2�񙸛U�/��^��ޝw�<kmN{�!����òؑ�<X/.�����,'+�B�P6�佺ƈ�������sm�@~5LL�ި���/>�5�	����a�Z�Ltlg����"����k�5*�R!�����*oK)a��(��ߨ8��F�����7{;ڽ��s��I��m�֚�XݹO�uwv���~N(hμ>k��+5d�[�͋��,˫�����!Z�f�RK�����H��J�ӣqVvȗ|��ɦ���Y
���1��yʭ����hH_�>V[�<P7���a1��a�����.wIN�����'e�T�N1"�<�&�Gz�Zc�=��6��Rm�N~��,-}t�M�ҙSt|].�5������=�I�7�!��:;;nWD6b��n��gh�c��3����3�W��lCms{!r7�Y)Ũ��mZ��n�d:�������a���Y��>��풹�ϪvQ~zaG��^�!qe�[���O�uy?�2�� �?�8tx�E�+��xK� ;)q޻��GhgX�ͫ���0��~��f>�WT���s��	z/,���[�߳}�v]���X�̟�0p�ZW񁏦Mχ�Q��}�n�B���|��K�f@|��L^.�zά��Ҭs���*������yO����02��%�$R&F���
}*���F�q��2���lr/.T�;y ���:�Q͗�϶|��R��xRn?749_��+;�Rϒ��A=��1w���.����)4،���8��fC��r.�uи��$JX-"��oKY�mn���{�=��A�qͅn��"ԙ��l��*i��:��D�4������Q�5ߍi������n���h[�@��O��Δ}wĖm�`_m��f����V`h�������C�����w8�n|̽J���.6-����y?L�8�m�?3e�9g�H>u��|�H���R�~�{���4��18p��dC����V(,��-32�xZ���p����o�2���IB�I���庂�+�:�4�OPO�
�Ŕ&�>pV���*�L�FyZ-g�Vg���F4�"uTD��觳���ԥ^i��M1��<�d�,u$o�g����Gh�_ ��7ܭ���Y��8�0Ezܾ8o��)���b�W��}�k�j{�L����H��ݨ�{�Q�kˇąuII���
���[���Wδ�5B���G)V
���O�fs� �2��[���m�@<����u�DK.Y�����&j�s��=��d(.�/�yA��.��V�X�Ϙ����+j��]vv~UȜϫ�0�D�{����p�������
*�=,F
�'p�X�I7�9�A��^�R�P��y�f��vך��Tp�u:�Ή'=]s	�T�Uߢך~]1�F��5�Ԛ�tC��l��/�߄�+FL��~Մ&�3�3�IM�y�*��V<�[J�$Pa�Í2MW��j�����Q®=��R�	��1��_Y&";T*ag���Ψ�4����㠒�eq��?E�V
憝&�%�x���Jx�,��"gv>��-�=>��[M�zHw(�V�\8��q�ҽp� �i2�����.U��<i�%7� �y����=GM��3�.��MA6�F���H1u�b�z��W��a��r�FT��9s�w��z�X9�A��������j`f��M�؈��
SuY���l��!�܆V��wLl�2ڙ�c6ɓ�9�̹�6@��*�L���Βk�z�=��:���n\��a�<٭:*]�<�G�[0�*����S�R'�:�^�����2��㊾�����l5�/��N�y�X�.�0�v��x��=���V֣��zkL��=��ъ:�W����D�&�S,��4Do��Fz��n�r�	�ӡ^�ae�63��qyH+�~�$!��9��j2&|��-%�x�So��J���v��,���*��s�� ��T��w�)>Յ�9��#:��a�fS�j���:�S����7ɎH�ڡun{�����R��`��7<��d�R^u�����9����~��P��\NY���M<,��l �%4�#1�5���L�=��>,�T��+�[݆���<�{(&�^.=�+1����s�ݨ�*)���;ߚ��T���q�R��!c�rI���I�<ϟo߈-
��,��	��"v��j
!u���!��n&��<��/�W��>�څ�PK(yY?�p�v98K��s:��Tc0vI� �(�0�ô���o�P������m�+����/5�Ա�>c�^���������&������\o���d�|kQ^d.Z�X����}�u!�2�؀�,��܉�Z ��V��=�/R|��F��hc��R��d��Ѭ��Ng�!�Jj3��[�%vp�Q7\�A1��9�������W�K����f�uF%e�.*�$�����I�\*)Yeٔh.7K���(dGM�ΜK��)�\K;�â�0��ץ�e\��Y�xK�]���;�e���q����%�x4Vm F��n����/��$T�w/��1����r� ��"*��i�\*���#3��)�^8�J�F������G�_�l�:%��hE� ��&R
ȥ��~Z�P���f�Y��S�%גU*#ZW�9]T*�5m
c�����2����˖�Gvg�y+adL�e׏��T��2"��g�$J�~���1<�q���A1]Dep�j��"L�J����}�t&6�Z�<�}���H��.��~�n���#�;�eP�����+�u��#p�&����3�_���r�}�M1E���6"����c����Dy���YX��2�G�W����R�(/�?���0��j��Fwp��.�����n�������ƈ]�('��8޶%�h,��$�>�a1�c���E�_�-H�/T�,��Z�Zp7�.��nPW�BZȐ}��Sp��]g�h���1f�lCm���ѯ�<����Z���!��3JGz�Z.g�D6IX��o/��/��kf.���^�q�C���g�E�%u�g��);eNx�>�E�̠�������[��$8����!fĪ�l�u�zDt���VMqbYX(Z���Ä ?�%�r��}��CT
��Ɣ_Pv-O���|�i;5��პ��:ūJ������r_o��-;���.�؏�h_��xI�c ��ٚ�;_[�<��b��ݲ�"VyCz��5ake|~����p0{�O;��&�(/�g8��'����O����U麐�r�V^e71����w�jI6��Z������}U9���i�7�t�=���H��`�l�\�}ww�Z�I�'`�x�o'�٨�.q��#�;�q��#ŶO1�h�~yd�*m��Q?�6�5�i��u�:k���q��S�ѿt0'��A��i50_��J4�T�LݹshuWMpn����F�(�?����0����GC=sઃw�a����@�h{���k	/�tE��[V�P��Q����0��\e{����t^�e�Ѧ�p�R�\z\vo��� 1@p�n$���x\����e�˻��l Ā����A�i��D2J��]��#�} ��+ϥ�Vv��h-YSTI�h]���e;;����ߤ���.�9�ת����T��H����@�(�A���,= ������>�`:�5�9'/��J����y�sg�0w�586�g0�@�u3�'�t�����DO���Hk��kw7�� ���?YG���(�ue�P�Î5ߨS/��Q�1��e���]�-���%��`���j��Mc�f�s������.��*Z#��9�����֑ ��xvz]�i���)��[������h�S�+x�w���&}[�T��0�!дylurH)��"6/��A�U0��/�W���[�)�,��H {o�e���q� h'���1$AV����V	O��C�H� ��Σ����]@9V��g}�Y��x{鱭i�(��I�-���X�x��~�5-,��)�V�"���5�a�ZFj^�}�)Q��e@e�*�5׏�q^k"Rp{^[g���x� 3�ο&�������M�o�*��:��p��^�t����\lj�w黍۵����g��z����Gbp����H.Յ�l֥�K�4*g����yuQ%Q;H�y{�FA�K�T)��.�7�k�g�|[<�/+���;\	5�)"i��.Ԣ��L�p23��|�ǃ��콸S�����ގ�Rj�e����\ʦ���>��
S�|�&t-�^��aIbY�+_���	6fh��u�h�ˈi��~�\�E�5�V�.g(��)�������GcaO�^a�g��1�t�����F%��κCP�\O�?{��&o3Z(�w���e*�H��Au"�c�<�T<Z���%w+�3�?���MJ�6%��]���\�x�����i]-9�{�{z/�w-��S��؈p/�dM��/�h����uV���e�����@�[R����.��2m_V�������.=
B�oe�'�p�������(<��u����o��	�Lq�f}s�p�Cr�}`�f_�,V�$\�|��@����f6N�.�s�d�=�u��֠����s�N��ĵ1��Z���p��ý�6�X������TEu8��?�;X� ������U�7^����luU�B<@�lS��l�@p�k�/8�6S>�ٲˬ��u�{�{a�n{_�ڢ>��Z!v>ؓOqݾ^��K;>&�#z�	�J`~Ȣ�pVf�/�}f��f��$
����(�/47N}���,��=�nR[7}� P-�u|v~�����1Si�Y���=R�����͌3�g���5�U���8�����E���g�(��M� 0��+7�i���_^���s���]��᪼-�D!W��3����<*%b�����F#�,�Qp�P�'���eO�8.�����cjs�Km�eώ�/�=���4��ma�qN���Tkv�X�x?^ڟ�fe�(�!����*��FvrgCIġ�%�u����%�((���5V&_m��)�4+�SArx�����L�\��N�ѷ�d斍�b���y��<�[O��a�yU-�+COr��� 6<ݮ<@�tSLY9�+vĞ)]}�+@��"t�ӿ�rԣx*��2�\İ?��_ES�v?�e���Y������L˖.��IYi7N�G�B��\6���po��Wtg=ö��D!偖�T�A��o�t�$v����`� �O3���V�<rn<U���UJ�џ�?�}C�7��D	��ҨU2&�p�*ؕJW��2�*�g�ϕnO��
0��Ǝ�9�#�k�n�0���_m��p�OcG��<��	��3c;�)ߨ?��>j�����C�5�|��[��6|A���N�@.�D|ń��o<��V��X��/~�,%�p����b�j}n����F�N�e����i��B�xsX|ր�f�2�@�މ׼��H���-����Gx�۱�2�h�����t��ݲ,d���������ٍ��[����"����%a��`H8��]��ء#��@��Ȯ5��y�bF~�z|��f�ö�|��g���N��B��'?l[YU,�-k]���޲�{�>"=�i/�X��\y<���1��rt����tEF��tU����j��̫w��KC=�>#|W�Y�� �e�j��\JZ�O[ȕ�'�Tg���{q:M��975���B��8\^��-O{��wp@�|��Y���<��L�c�7��t�g��Զ?e��2���(�:'ѣ�?�Ԛ��ћ�v�y�ԛ�g���c��P������_��9pht@%R��~/��XK������aB=?��`�M̘��p��������1� �1L��$#��B��:T5��~\��G�F*�E���7���s �:/m���{�|dM�P��&��YhЎje�$y�&g��)���@8)�����bmQA�7j}�9�ǤZ,E�(�pkh��VHQ�Pk$���zJǕVn"�Uly�� L��gϴ�o{���43l�r�C*��4��4_���Pq�:%��PJI��7y�.�NucV/j�Q�g<�ft��MML$�i	�N�$���`��d��5��}�.���p�i}�-!Q��t a@sG�nSV��&�E��m���Ty�&�Z��ZWH�_r�����L��q@�U����b�6��6a��\HHT|aƪN�YƇ�8��'Ǆ
������mƲИ�_��2��Ekq\k��:���l������M��� �����Ч��!�Րύ���d����*��6���������o��|�>��S >�^��:�S�*2��{�ds#���"��7CL��ݒR��uS`b�xX�������c�)���e1N�!�9l|��g.SM�2����(��D)��>�O��`3�-Gl�=��K1Z͑?oDf?Q�I)�OL�c1��g��'[�< QAT��l�R�2`B������Y��0�˔#��m�� K�Ailb�{��}R�&!�b��vmPt�c���@	u0K��Ȝ/G٥��xK�:���!\Ut���x��Rn��ze�/8$��e�Oك�LsKl[��H����[2��G�x�Ҏ���aG��B;�&/���D�����W�wB,߮6>�5��r��!��~;�ۘ$]��������I�[J��"݅Gk�;¦\�K$��Sve�M��مuܙ��.p�e�A�a�m����8�QI���z��Zw�cI���M��Y6�;�����f�z�n`���筝�V��������o��.�TD �=�V�t�������;l�.>Ԡ�!��Xu�S���[�V�Yй$.V��G63�~�L�k5��ǭ�ȥ�����2���v	�/<��R&\k���	/_=K�gc~��H��/^(���G�׶�M�+_�ͰU��&��='f���.�HMK8aeC�-��t`9��r�t�c�c��������H�����2BEE��\ΘUq�H#���qEeBMyQ�Q�B^���u2�l�D*%f[���e�W�ė[����ބ��w�^ ������� �Qؽ\�yIOxY��W�@P �H�8�q�;�3��G�7���*=�5	@�l�Pg4����8ރ�d1e�IIM��zs=K�h��!0޻��P��x���4���+D=��=�G0c��4�r֭���3ml/����i���㯹n��n ~�1uݡS-OQe1MS/��Q���s1΀1�5�9���!� C�9V�Jh���G?G'��BR0;{�B�����Yp��n�c�%Bl���$��ᣤ���	< ��ܻ'�[�`�o} L$�hk|rHt�����=I-��\�~E�S��l�ߞ��@){vm�y�F�U�6��@�W��ɇ��պ��"	/ 8895�i&��S`HD��v������@��T�
�Ƴ�{�:��khi�1Ӽ��|����>\T��,�z�䮅)<�Q�@�@W���k���ܭ��z��n^�o��C`{*���xS,��軑��Z�a}�����P`V���µj�Jb�:V���	���;�(z
���`�[0~(�.��`�eQ}W^�X��kp=�'<��>i��_�rL�J���(�0�?���*^����\��b�`�/,�=����os��"<D�ތ癣ݭ����Z��Q��`�2�}mu5�a��P�X�	��RV��
i�ͪ6:|���8��1�Q2V��QW�'Mɼ��r�Z�OZ)=s�W��R��#h@�m:ѫ��j���<�� z�A/[����<����믅--�i�!��hvRRrb���K�M�.�T��� +�7��A���������q`-���)�n��*+�=r�m��꟪U1��i��hw���7�U���a;!1��'DO���E��*o�B�RT��������̏ �(����d�H�K.�ߖ��O.,��8ߎ��U�W2V933�	�	�-6���ϓ�)��(�kߔ/�n�ųHSgI{�ǉ�������˃//p��(^O�`m�t�ɿ�|��ΰ5���傔��3&G�_�E�\�G]<�}�=l3���>h�zF�����_�ȥG=�D=Ѽ�IF:��ຏ�i�UdJ%xz��W�����9�Dv���t��в'ɒ�����7�=��j�|T�op�D/�"���)q��-t�{Upѫ��;#��q�삑���RA�Hhr/|� ���`џ�7`�,�.���WJ���`�υR��;r������Q�����AXm�\�b0�S0������9��a���b^
%��."�:��	��r�C�	rD���ꝸ<����#�Ǯ��fGzerEOF�v(�$Œ��U��f_�q��sB�u�-�.O��/&?8:��E��BMIX��H'�e�|�]����Ħ�/H�S�٧��V�l�/��y5�sq��j�he��݌/��y��Iӕeo� ����1���gk[F���c���q�2��9��K�̅4N�ݭ�ƪ,�M�.�M��b5��/%A�y,��wGV�{,�GКD��-�&-M�.��n<��hv2��\|XX��Z�A����9-bxxx	<E\5� �ڲ�OD�^ť'��Ȧ���"p��x[�[���˲ӭz�C܃:�ٵHх��^�<���0+�56�E/�D��Ũ��8���*`0 ��̃i���ϰ���bb�+&�:�Y�U���LMMkڙ
E_��'�Ƿ�0���Ɣj��W#|����(�
N��A�=-�e�A��>>=�N>0>���H����v�V��	��0Z�$*�|��f�ZYY!N��w�	u�X�."|%�YZG5�F�hG>-T�Q��uwu��V�}�J���;���م߼�h����өY�9�*='?�V��%P(T�ULJ
<P�:11�[�_���?��0^��>�k��6RY��	���y��y��G�x������u$�7��kqU�p�ş0J�2<�^�nh�	;zӐ���=�n����.P��TǷoy���7!����d�k�]g�`��B��d���Z�qh��X^�� ��'�b1Ñ��a|$��lCԝԟ�OM�?;�\1_�b���j^7jd�N�y �-���x�A��M�d�zhϡ�9Ɵ��ADh�k�CZ�hj�v�Z��χ��q�=
,����������L�2˃XyM�8(G �eB�ج�o|��8謼���w�kz�����[7-�3�%�r�s�l�KP��_m6�ub>o7�
��#�Z�7hU��<�'D*R��]ID-����]��B�6%	�iw��}۲��� nn�&����f��D�������e�\j�ty��[�Φ)�ܪ�:�,�}��L�P����zY�c�ɥ.z�P�H�����x�#�������}=-44>��_FDn�6N��ʹ8Vv���� V8,��H��J.� ���|�g�5ӬH���mJ�WX�}��6̸�aFk��}�o��FE���H�B��Qsp�[��h[���e<骎!!�%��v���n�g�qjמ���/|� 'i�#��8��nG�`S[/]�E�$��']^��Lzw˥���z!ºa2W!;����~G��O=�����?}@��	Y�27\<�%¢Rv���e0�9��B�]��\����.ZLwE�c�D'��B�8F�}��{�F��g��Jey��Y����l��}GV��uq�'�G����PݕOW��:����G����R��T��=��kG�$�&&JZ{.v*${�{I��S�ӄ2'/�NWRSJ��;�A�g���ݨ-�����y�y���g���
%��R�@����U��z�f�9�����#j:����e㌲������9>i���7�z�=���_��p毒E������f�T��w���a�G5������CN��D=�����g����f���_��}yX���1!�95�3o���_�b'<MWfh'��-�y/�ԴC����af��s���R���>׫�x;�>(,�u7<P�д�1��[:!!�݉苎��/��۪��4mu��l�I���)�}xϤ�۸�.��d�Yt���td`#W���Q*k��X"�`�J������M�d*#uK>����rb�3&* ���)v(���fW�݆�����=WiIt��w18� �`OS�J(V����$�,11Q� �����&�fACv�|���p����l�~��Q��@C#����s64�Pr�������{l�s˔[ �����ZxΈ��L�ݦ�$��h������|g��ǒ��@:q�����n������}��#����=�UV�� ���Y󈉿J��8���$�����4�H�	�hD��v
�/�^;\ }X��N����\7�z�����<P��`���Y�
���iH�98��[O�ݾo;1��	\)Ml	��sp�[Òz�\�'Xt��#җ%S�b����6f�>��uu�tŦ�ݶ����mW{qo=�༴��2h�׷<��&�S�;:4eh	1�*ߪ﹌��\��lͺ��)z��0�w;�Vm$ ���Q3�p�ƥ��o�1����9�����K�c����Q�v��2%Ie�tl7���\���B7 ��a�?�!�a������ٖ�P��8����|�
���1=ey��#�%��O�p���)^f�+L�
��t��.�� ���
p].�L��f�{0�ż��@[�`���(DN%'>�;ʵ�?��.���LBЄ�����C|�t� ���H8���-l���x�B���s����>�)CS�O��#P�y䢧ݨɻ�'"��3��� $�|MHXrn��ˢw\��!Q�=2E��7%e�z�q�jr~�g��.���a�����Z����>���:D옟@_�n`OJO��z��	eD��A6�9�*C1�o���G��W��3�w������U�G�^���)f⤭�<�\xǦ�[��B��^pD����7�k�!b�/KA�_�^m��1y~x���KF�-�g��ٍ��������Є���I$Ȩ��P+�q��S��D�m���h�Ք�@ ��\��{0�Ii�Y)��sTx<�l�A��DS�g�}�o��~~hHy����/�(N�0��x�0�O{���9���@&s��i�H��I���)b#3�M�/�����w�}�D5�8k��z����u=%�u;��o}��%vrŢk��7/������_�y���Jּ�b���(.4���l�(��U���6�~��4�'�E�|}���d|��X�R7��lD�׊�nO�ybY���vBd'��mB�@ߔ"V�-sel�Zk*S[��h.IG���ąc�KT3ڴ�Q��jWrB4�c5*�N���o��I�D�>��״�?\����V���
�h�M�r�)�8����Ѣ��Ngۘ�$��$�PK�n?���C}��7@�^XL���
�=_�Zp��P�hA#N3��@<���9E{#C��I�"����v8���9�UD��<j�EeX��=����yl��L�~�z�7ڬ@���A����4�i7;�6VO?��7P=�� ��zB���5�m՘g�)M���|�l�շ��L 2������ax�V����>��>}J~�/��J"��#/"_[���@�� ~�rk��K���i���iưe:��?��X�`T)���Hm���s��; �k���!Oc(�����zb���+ybl�?��'4:tc(�s?��ٚ�|��cv���H�~������\�kg��Mڮ3	��>Ҿ�~��kKI�E��.�M��@Ko�e{�Jj2� �վ0�P�?Sd�+[FS�͡ՙu�a�!?���7(Ȓ8������K��x[^��o�o=u]?R�������V����U+�a��3�gJ��D�]5��GS3jF7�`lf���uH�Q���K*x�
C~]O�܅]�z��F�kp�ff�?�b�F��
� 7E|�7��1�@�	�C՚�q2vU�F���<�U�t���a��Ǆ��s����2ɀ����2��7��]�!�+o����S㍉� �''�<��k�_��U�%�`~��cgSŗG�0�/�u�t�3p��49m㊿"T�9����2�q��Κ�}��T���e�C��N�Qr6�nM��<w��eLp��z��
��I���{8��l}z ���3	�n�(�1@���3�u�[s�~I���􌱦�)�L�����@��ܴ�|�Y{��|}}�����5d3K�u�7�����/G1��5��@��_��5���^ღ�W��+C���Su�Zz;9n}y����:�W����8C��;�n�?�u����������d_G���Y��������w�k�w��V���wH�Y�Z�#g��;�*�L ߣ^����l�O�D4ey٩߉D�����В��%[��BsV�뚬 �q'��C�(��_����g�bʟO�q(�^okl��C>��4ט��x1l��^7u�vwݤ�C�;�Y����I���p/��4�@T1·]]��}6P��[�1�z�ű6}gT��Br���j=}�B���M�Ok>�_<���O���%%%)��LE��7�G����ݺ�ļV"�y�O����6wv���-�m��hXk-M�B�������ML��Jl��$v��<;F���Ӈ�,��bs��}�D6?*я�jI��Ե�RYI�/��� ���u���d��xe�X��e�;Q0������-�^	E���;���:���5��ıWYf�J]�M9V�\L�L%�������?Z^�O�_�q��ʗ
n�\V�������s��]W��.�ض�i���8�N�9m�>�������I ��Q(�x�y�s��t>���t����K��� S+x8x���u���o������X;E��1����h�Y�$�ϭ];��>�	@�C����EӺ�֙wh���.�]���T��B�V�H�i�����H��wO�ۗ� x� ���n���w�&�<y!��c��)Z��x�q �S�x�2��_u�-��iwX���27H��$ ���\q%�U�xۑV���8�t�%�10�E*Đ1����J�6G㵤gn���6��B����� >�=;�
�N�)�Fه[p��!�V��V�tL�{�kGW�/f��{rc+°�C'++Y�`� �8�����?�Fp�)�d��#,f����������8IKK�ى�

�f��9�+�G6���4`����Ht`
��d�Ϛ����E	JJ֚�����Tz�6�Ԓ:L�����{ ts����=[t��{�U11�D;��J-�C��t�!'�}n=G��)ˋt�㶑�8�:�S���^w�\;\{���V(z5�
=�@�\�#e� 47�C�Rb$� rc�7g����F�ͦt8fN��u_>�"��yQp�x��Ծ�mӖY"Yg$���n�\�<�'*Z������P"�`N�,��F穲��5��#ז�����D�kh��WoW��몖����o3pi���M�?^�W�08O C�ı�ݵ�q��췇�M^�;f���{���d���a]nݧv�^b��o��UF��BEGI)���b���4� ϰkS��ݲ߃G%*U�G�
��Tj5�t��zJ�ޔ���z�$~zL� v� 55j@�4�t75�^?�9ܲ�j�.��ދ���0e8�K8�p���%�;~N�p��Uw5���r��p�ȿ�|{��\JUT��5�K�Ąu��wBC�^g����fU���.R�i�_�N�^4��O������͗��k�l�Sq�V����i[�_�7z������z���w*���+MdG�gO_u�b%�<�꺱N��F�螣G�@P i+��@I�1%y�=H�������Z�7�2L�.��2��g���n�T=,t�-!f?)3�uY�t�R�9���ԝ۞��8 �a%@B]Nc����h
�g`���J;�Qnnl���/T�&��4�e|�;�+��2A�w|�q���i�Y-+-� hkر[z�:��I�9LU맔κuh�\�Y
��t�����V�E���>Mڟ�y*�^�/�h��׼�p�}�ۀ����ŵ������ͻ]��������R�?)(�����+2I���O- z�(���iMXZz}]�����~š���&4�H\0��CUM[�C[�����=�`�/i������������2�_��Z���7�7qڧBi�ox�O/1����>�uW����wo�il�}J�X�{y5X��M1��������~[��d��MIOQ�ǥ%�L�Ώ�ф|? \�"��qV`c��OVC	�sQ�ǗkQ�;q �Ŏ1_�[�:�GNn��ϟ�3����$ Q�s�?`E%�)൮#��MRw>K�Ի�K����5U�!�OK�J#�Ȫ+�a��Q��#� �w��m��+���/oX*��2
��O�.}
qt��L���\�E���X`�o�i��������QQ�_��H���� �݈ H7H�tw�4�-=H��R�]24Hw�=�����X��5Xp���|���{i�;���c�.��n���,Ro�J�fk-��J�m_G�8P:�+�k��0
��z�D���cn	�z[q`ٽ��tH�����ڔ��/t�{0�,�=�Ck ��n�H>������:��ѻ��w��7ʪ��'����h���e7�tyqO�C׼p]�v2��R�y����������511����$�ˈ�i���ƻw���,�|��,<=S�I�|�������N���3Hm��6���}i� ������G�W=$\2$x�#��J`{��N:ۃgX�>��HY�׀ԟh��WYë�hP���j�!��<�m}ML�e��gy���*�z�]�;O�M�!Ȫ���Ի�yf�l�	���,��9]s��ۓ�X�-�Ow�jV����}�y�U��D0Qe���8n܊L�\~C���?� v������6"�	pa���������?�3���X8�O$R!E���V%M��;3�7�_�k%�p�.�﫯�K�'ةUe���~��q���b�z7X�J�VU9~>��x<�\��\�L�ч
��h�ri@����a������pY������ZU�0��sK�A�=�����Ő�H T��! ����� *�-����OOmmЯ�ƺ�Sv����V��|�����uR�k���m�4�b�!9EDY���J�(�z���S3@1�lK��E9.�����];[69�����p��Bm�����r���Ђ~f��;%\��Es�OF�A�����b�,SL�i=�i���eqs_���(��g���(���Fb��3�=X��O�LYC!���lOP��Z��83��l�2�8Q:i4���2����<a��VO���.����&+���"s�N\
UG�S��݋wR�m����㬭jj�y����+���\�*�Se]��A/H�r������ĺG�B	d�A8��c21YGxn����P��Sl#�px��5�/8�ٔk;TH����������]��:��Ǜ¤�16ğ��4��W���E��vaT���B���j��H�>����=|��jjv���#I��Q+�n\�j�TWm�4J�+���?U1lL�d��.? ��j���	��o1%0^e�u�����o�>��b�H.�ߓ��=�6N�� � �Ι�ݯY��Ϯ��q�ekN3*��a1_��KMÃ��LS���*��dBv��p�n'������5��`�2_����B�[��y�ns���v���ߢV���e�D���~�����&����d����>y���q�� 1�g��ƸV��tQV���:����n�Z$s�s�k.gb�^�[�h�5���f�n��o�W�)�:D�T�o��l{��n\�z�&�眪��Sĺϱ��3���s3w��㚿�%4g��]�=X����|�t�j��5��`�PQ�͉�Ԃ��Z�¡�b'+NΟ[��uC��'r�c*l�		��M����
)�����J����US�	�dZs�c��^<��c~gyh:K�J52��dԐ�д�����V�pv	$bpP��� ��pƗ2l\Q�����+�L3 ~RǏ��h��t4��Ŧ]O�lQAC�,�16U����K"�?�ų�yb�۾�n����YD�6Ɖ���;���A<�_4�J�2����O�]���-X���c��R�Z��/R�Az��lߌ3��������4B<��3�;}��4R���T�ux��5�"�'*#^O�g�7B��׆�/z�>�������@4�p�@~�8l�L�)2�q�DE�Ţ��'ϡW��U�|F�UQ�oP���ob�S���c]���ը��m�X\��Ax���'�?*��f{>�\��;�t��Yƾ�����$����!��]1P��3l�Bz�&$$?�ۙ�}U�$Ϝ�r�r_Ub�C6�'"eS��T�T�id+���w//���_zm������/��Z���v�j/��Ч�C�(5�5��yƦ��UoN�5Ky�]5n.N�mOw	�������6Aq���s����
�mE��5��G�>e\���Y	Fe	�w�%��`�����7��iD�|�\���>����*�A
��-���G��O��B ��@W���9�o�'t<;�E�:I���q^�4�.����w�1bQ��9
� SX��{�/�F�s�"�&��������qr]�+Wttt;oN�N�ZX�8e��C�ɨ+F�w�f�0�qk�Ӳ�1f��^��e�% ���WK����o����F���	� �9QҩS��9�;o!ӿh'\<�$j���ג�:;��5�>��_��s?���̆#���ߠ����G����"Shf0�ve�^���S�Y+�*4s=�0{B��dD��_�(�T4�PĐ�YurJJ�����BLL�
n���
&h��.F���rIF�jt��=�C�ʾ4��:����Ҥ���C��ސ��;'�c�p��]��R"RR߾�!�j��	���Y푩u�X�G{����{�,J���hk���.���������8��֖o��\��
��+������QZrϣm�^<?l'�0��Q���n%s��!"W�"��M����Gc��Y���{WBֽ�&
0�J��ތH�2\��`�X��n�[ėR"��|Q �P�H(��7ˢ2D^T�\W3��/�}����-)r5��2>~	s[�Xӿ31����p����z��>(����6����v-5�tA�V��G��("a�G���t�G�K	g��%$��E��=K@��{���TTt�+��!�VFg��1>;�.N
E�T
�K7�=��q&b
�l�u�"��}��>#{�<Z57!����н���t�Jw��ۖ������U�'n�il�ET�� �������Ky��~^�����ϒd>x"w�1�n�z;s�� V��"��"�5�J��i(�q�ˁE���/�Q���K�_��K*(`�2�44�#{��w�����u��S��_�vz��ccc2w��b��a���"��I����/&=��'�5�]���:���
VJ�o�"�Wn.�/:Dn:L��+?kNp9"gH	;�!��)+�)�2��w}�I~fS�թ�A�����s~�ޙ���J��#����FB�OE�����9�_8K�^�9�޳���\z��sً�&X��ћ`	@"��������Y��#��
���[9q��&�u�Rd�_'M��c�;��4ajj
{|��ѡ�h�Kc�ڀ<Gv�.�Z�>v!��B���|xl�ӑ�l�".���	�t�%S�;eJ���ĜI���NQ��K�+�ٮ�z'ۤ���o��)�}�/:c�U��ĄC����uCƻXt��"�y=�w_ J����v}���~����Z/�AdNgˑ�[K[,'ҏ�w��~���\�� ��C�6�7����^���M��ԡ���iHL�b,�\I����K̟�q�"ݮ�7��=�b�v�D�0 �GҎ.��V\_�{�͘U���R� >?���$Q<�<�G�7��8l����ˋ��\�>��Ҏ�+��y��)<�H
�:\}��F*ɹ���uJ3F��9v���F�֪~~��s��g����C�:\���>JK)4����q0<:�n�eʀ���L�#��j�A��E�B��L�mR1�a�S�wT��{����ɚ��Z}�z�@��c�X�pJ�V��ML���r�VDU�.)i�h������^�������׭O����B���\��1"��R$N�J_���ȊEGw�_M	�u�ϛGh��.��E�b"ަ�;�y*���"]��!��ၛ����ʈ�O������;���6i����OTp���@��5��y���N��?ے��k�	�)N;;y��D�,�5z;��^U��N��_�M�Et����q��i��|��e?5LEN�c.��_fF�5
i�0e,��)��BTD$C]�a�l:x�ͧ
3�X.k�#��	,���D�c�첅'������"�Ps��{�}�ފ�nӋ	#A�5�Q�m⓬�3�D�i��J� �!�G�w����6��x����|��^9�h�~.�=�������KӏÛ���2����Dz��w�r����Gk�G� �����0&���+�0��.�l���I��s�FNV1����`U��h�����p��M�B����@���V΋���f|f�o���?Ǆ.γ�n��2�y��OuU�ڳ}&ː3d�E`	}^��ó�}r�>N'�7؍���x��]�l�}@��7��I�lez��i�f:\ѯNk|8�O&%]�PL%�$��Nj���®F��
�w��.�~ɉ6+�����\1f�c��]��\+�˰`����l�̢7c(A�4^��n�i�~=�01I:5Xe�$�ڦR��~�C��݊%n�d$�ٸ$c����U�.����o���Om�0y��~�Y[�ȋp�4B��a?��Y�?�z��~�n��?�}���弯/�60F�sI�O���E���/~��o�{	��`ϻ���^�ę5�@����	Cb���CE�]?>E=d��c\P�hr^��������/�b6,W+0_
_��{��'�<�e����U�?�mʦc�/��9�p���uzk�˥�2�«�����*���"�qY���Ƚ(�+g{��6�ܿW�9>"�5��+d���~zU�'�#4TȆ�\$|<��G�M��|g�P�����2��czD~���1�W�(���]�����3�J`m���2D�����S�scp�D��2�& ڡ���k��������
�E.zx����s�5s�f����v-'���W�c�g�-���v��a�A
ގ�w���kA�
5��Dl��7W��w筧'��7w��V��=>����{��#n0-z���[|x��𘅸��\���c��ӋlE��-|9,!��G�
�X��+Gهm��\)9�>��@��z��Z�6��H}U�o��_DtR2�9�^*Ȯ�g�Ǽ�@a�\��z���#�c:����A��N��� W��h�)�����r�h�RS+_��U�Uj��:2j�d�/��4��a3����:l>q����
xB�G׏/�c �_�ίs,&�VX1���f�	Rd����5���;ׄ�q*/G����Z���h�B�l6, ��'�5�H|D�U���R{����5Ƞ�����u6�qC�Ƽ�窢���������+�q4g����(�Vjb���5��ev����?4�:A:G���悼	�����w.���棍T�~���q��1~\"2R �/�~�5�Ԝ0lz�y��G� m��K�i� w�K��^.�AJx��#Q��]��'��%�+צ1?CbE4wx}+�&>��HQ�-��o�89#�sgǺ3WD�#B���U/�SY*B��-�*���!B�}�:ZC��%*�W)*��z����䴴^m9c鋝���:����A|�n\8]�7��qZٳ��_؋̏h�T�%& �E�rp7�(�"X�1>�*�Z$��R���#YɨB�ƥ�)��c+�tZ����_5^;����f6k�����܌��H��>�^�::k������'ZkST̖�	t���<�hqb8@WW5�d!K���lH� �7-��r���'T��z�����r+9M0~)�
:h�>[�G������{�J���TIWW������2\$-����B˯�ηߞ�/�6�%��󅉡�ll.��p��׏s�˱���.'���m����#��'��A�HY,���.�]�P��Ȟ�0)nlF��ٓZ|7�l���#h�t��uk^��aP���)\z��XO��,����yv��׫~�Z�h�H�����v]�F\>�嶛�b>^�zj�����A_"3��"��`|lj�'��@\�x'mK
��a�o����Tgg2+�@6������1��łW��5w�XЋ�X�Mܤ.xT`��l:r�utE���v[+���[�{c�uo���������KՌ�׏U�ʦ(RR-���X���d��_C�'ss����>�,׷D��bff4�_��"���l�oT��eoi5�����&�]�����6F�&��C8��(�D�S~r$	���������]�A/��X����G�zu����D�2R��J�c��kw5iԀ��h�j5��W�o0}�ND�ד���U�������W�̇i2Bw"w]�PH��B`c�MU7Y��4� E2TI##���+�7VO���X�:u�)h=����鮪������2�/5}c��*;�X5��ev��as��/-P�ְ��5�����;侓i[$c\�urv�\�פ����2޻��As��{���9	� 0r;���:���D����iY?~�w Ʀ�N�¢�u�<�j�H�'�lCՖ�����g��|��ࠧ�?4	%VVV{9�����L&%r�e�8��H#�v��R�-�S���g��d38��ߖ��8qCmS
�ݥܔi�1{xYY�g�dM�����s�J������(�Q�����z=V
�"�ok}�[!��_C������t|y���3��N�b��"�adg*��.֦���궻�'D鑹�=e��D8�^��状������_S�;��e	�wգ�H�}Yi��@�6�<�������*�./��6 ^־�Pe�Ƙ����At�S?� ��7���*�!�y5=[�F�\T_?l�a�QJ��
#6�����pu]t�/��)��(�1hZ*�sg�˩@SM���S�yjH@ \: V�INcg��_ޯ}�%~.'��x���v1�_�f���.|�פ]�lw�.��>�����?�H�W=�����X���~%�Y��W�gb6e+'J��P]天{)۾������#\3]h?b���K/�X�5�l������Lu#:�H�:��W��ل��m�����Ϣ��k���﷪Dx8g7�O��x�
7'�3�:W��`JD�dݕ�(0f�F�f�����hc7��G"9ش�JW���?��#���?3Q��ظt|	��{���a��#��H� QfF:�w6���o��6Z�rE�*P|�o� 3iLn>ЖF1���%1@tF_�RƓ��?й������'9qY�@�(<��:�����=��9�غQν�ڛ��5Zy� ^�`���_�b��v-�������W�j�ou�2�q��hf�s(����p��ʫ����}��h֧�f�zkgǂ'���I,�vv��w���x۝��Ү_ ���Ct���`�/>|�^��	�Wo߾@e)S$|�U��|��Ƴ�gE �[��5�/7f�;5����&!!�k7v��d���":#@�2B@�P��i��!�]WJoػ���9�%'Һ}��42��k�4;Q�6AJ�H��򾖩]6�RT/�]Hj�BAIU	�r�A�@�N��(Sd������P�]]�k2~�3���_��L-x����`5��q~���h���F����b��<���gg��aj}��"�B�M�ڂכm�2	Ȍ� �"O�m�M0�	�R>G5�.��z�w�L0<)=�䯨!�}����Ԍ��Ы��E������81�8��p�t� ���Zy�x0��w�8�Ԙ�qqh�g��M��]�K?�ڔ��V���5����|����{MM�Yfy�sx R}pN��Ki�|�ϖy�[�qjjj�?F� ��I�õ��6�G��]}{�)�?�����ʿ�"D�Z^����[�e`��l(#:j��1�ȼ��ڭ�+M#�/�ܹ���坑<����%�u���s��MHϐk���^ �K����禷4"kR"ᚅ~PG5�|q�ٵ:��h؁Kn�x`��׍&Y�9�L�'g_CH�:5L�4��2�e�xz�\�1��TX_�	wN�Ӎ���ߌ�E�t$�;��@ԡ�r-/��^�ϸ���z�8Y����T��5����{��e��ܭ ��F;;�-dK�V�̚�(��-�A�Vu?�
[a5c��fh�0��Fq��(���0�y/�_b�8%���~c)��E�]_q���g�}i/�l�y�$��� �ky�7�5�:j��k�!��"�H�הo]7˃)Ajc�'2%�Ǔ�3������+�1DE�|6���㚅&4Y;2�'�!�$�Z��0~r]�]�kDRΤ
��v�t��G�z"��<;9Ǧ��=2@���Ҵ���jE�KPH��6�K�uTw��D��%F[gR���%5���fa��~`G�=��r�����="Y<dھ��kV��Q�{�4}�r��"ML�����ҏ��pF_=�.0#��5Z]|E�� %?�c�1�����=�6T���]E]1��M�`h�)��t����;l��ݳ�4k�����0;&�w���Q�d����7-�[zܜs�3�1��MO$��<L�r1c��T�\u}�@����,��U{bgܹz(�\a����a"Z�s]����dh�b��[q`���X��W8�u���Ӈ~��Xx��Ժ��A�%t	��(�9�\��8��ޔ`�Z�D�a X���w+��""��G O/�JTJz�J��p_7HЋyבb���(���c���۽�cX?�Ci�ٳ��A�}7�oL���C�}﮲���',B���-�,���������'
.��a�J�[�-4�d����aA$54Ԩ�\�B�8He��tb����kr��U�;x�K�y4�}��e�Z�xy9l��!?$�t�$�$=Z��d��_۱j�c.n��0l�{B�����PR����B8����-w��C�c�w�?|�6It�\�n���#���:���|��(�3�b�Ю��wY[rսYUWR[��A�vu'�_M5-�|�;�gh�?�����yuf7Đ<!��0_�Ȟ[t�g�w�q�vrZ��#��!Q��m�YO~����ֱU��5{&��!������+�(#xA�Mw���8Q��`#�{8۔7�:�HR������Uｆ~�!�߸��w�e~����	�T{8ʗ�/�ł�x3�Vt�Nmi���ô���$$�(��/ϰ~Rǅ���/l%�F�|�T��tk��\�D_𘛳���c1��Z^hh��e�;/��H��j�����܏�֕�s��wW���w�[o2�K�ھ��tҎ�L�9�ϖi秋��{�����K-n��y�L���d�8��[���v������9��þ��!�c��*zI�Ym�nw�J�tuZ�?Er��~g�2�L���>�`��{����1[��0d�n�ϗ�W_y�Z��SE!�o���v�yTz$�?M�N�hV�$���U����8�-�������y�}�Dj�Rh�.����%���N}3�c~'�wr�8��2mY����������濲��O�J����^�6�*�>품�=��(����z���L� I��	���`dܣ��f��w�*���,�.o!6�(� w���;�f�r>>~�w����Ǜ�u:�P������pwe/�����_�䛱,�,��5��j��ɺ��x�pa_����T�$�1w���]���e�tr��U(��3vJ�&-Gę��� W��}�sњEV�5�p�i^��5��hnqm��l�K���ϧa3��{�lpim��l��LA	�H���v��jԿ^�DL�Ǝ�̰�b,е$��j8-��T݂�g����@J�%]����qMJ��;�/�{�2���H@�������C\�m�{�?\�G��P�B�}�_e��w8.�e�7~��`b@�4���o���P�}�i���XѬ�^w�}�j��L+��o^�\�
�G�s���(��H��퀐l>(L���Uw24������b��tĽ��K�_taPy���جLe	���b_s��?�a�߱'޿?��K�oЍx=��Kv�Ɓ��4��P�L﾿"�a�$�1X��^��M��Q^u�bVFS��t��n��1�[�vU��Κ�{,��=��yq������Ⴂ�|��	�5k�I���&3�4��~>��|]B`�l���8zS��j�����R,�Q �5�̧�B`����am2$q7��:cA�|�:&�g�9���F��6�KIoy���il�EI3�$�G�N�_�y_�������l�d��!�8��*C&���Ve͑v��U`15���Vc=��o'kQ]�zL�֢����<�	3p.�&t����Q�9�S����@r��P��{���w.JΡev� ������d͜��M��|O�v��x�&�h��ͮ.���	��֬Wɿ4�~8#��Hڌhu�}Y[�BҼ� rV�����u�K�.Q�7����Y��`\��I*��b?(?wJ�~J;�~�Xٸ���j�����O�3ow/o]I�7�Ԃ���Q�&S�O'`�
.Z����]�.鋴\���ؗ���`���n-��7un�H�XP?D��-P����v�ц0�)C|]Wdaq�o��p�S���j�;�� �}O������ɸ� {�njY��o�;Q��'�F)�_�Q����B�3�NK�6��G�wϦ����L���������q�E����l�i3�j�ژC�����c����l�瑟�C#迃@�����׳���-�m	%�0��1�~5Ta�Zñ��-�<��;��L�V1y�i U���e�g�"e`�8�o0g��Kbq+jl.��Y����7���pE��;���1��*�.��I�A��%�IZE�ngc�s����Ǥ?�D�ۜ�f7���5�4��S׬-!���t|���̀ϩ�yĹ��5[?���8G���Iş��]xyh�zY�cu}D�Jz��>b�Рv�'\UB#�q��8�`���Z��9ҟ<�׈��u�����-7r+�j����yoq^��l���Y��ۙ����E��SpH�%��+|ks6��� �8��X�4���W��s>��*�����.��n�O��8�ķf���H�[!�϶��NT�d���$�_��ƈ�T�}<쥅h���3�?�5�F��S���fw�� Kg١.s>�g'�si޳�La��7}Θ��� ��y����|�_LOG�x�{�9<JMVa�{$��jⷧd�igxyM�FŎwc�
i�߮�@�ީp��u��Ǆ��Fn
('_�a�9F�������P{��@���'l�YU}L�.��a�]�M�-��K��.�����I�-j���0Q@Gv��ז\r��䞞��p�h[�_�J{;��e����=%����l��Y^9�+	������O<p�s���h6�"�{u�����1�'�ô�G����}]����A�����?>5b���n�[t�~ϊ�������
���dcu����I�e�Ϩ�,n{��U=�'�I���F�E�ȿV��%v^�� �X��օ.�~8CH���|�������ˀ� d^V}� ���כ[#փ]
,)��:ߣ��6�aH��r�_&�����a�2���4�Kc���Hz9eJ>�}4�c�"���0Y*�7���{�n�MXq�9=�-@�VZQR���h�/�{�8D��0�,�uw�P�����Ѥ�)q):�|���ð���	Gyj蓇h��4y2��b𵮐h���I�B�������"�x/ݓa�������Z�k@��Z�G��	�3��k]��0�?�6no��3��l�2�hL=Tk�A]xMf��O�|>��u�Z�%�==\����L �۳H��y�e\u����V+��ǝWBf���^Iu�_�ʃS���J�qQ&�*.�E䁶W�tp
�I_�4yx긃��C������,ѩ�N����5M��9Q������������-��
�@���l���Fr�C_���>5jRR�����XU����阬k�{�ǶR�˓�ۗ��9}�R\���#��,_wʙR�`���;Ƿ�����0u�	�Kcxbx��¹��1����Z���wv���@�[����ġ����O>�T��\�K�=��av���S.�n��%e��P��W���,��S�s�f�B�Tm���N�޾j
Yh�!jk����y$;�o@;;��N{!���
\�u��Uڢ�9o1�T/������ZZ����V�ˁYtX����h&l���@<I7\)$�xʢ�^�vW���=�3����O�a`�w���H(6�����FK8 �C��������'��=���\�OhJ�4�FEq)ԝ/��޾柭\@�gSu�̘��'n,���٤h��W���,6����;�/dFA ���#�\k�혣D��.��U��Cc�5�ARW��Y�=��O�������/������-o���A���H��QNt��^��
��<V�*��a$ �K��ۺ=�X縷��>���v�����o���$	4�pQ�sc�[��qw���ߌ��-�Kj�.���˧�̩Ӛ��B~�2/P��ʗg��!����!}�Ãl�w�j���'�K�=)囜C<���WFng�`.��˃����%��u�ձ?�_�����F���ξX���̝��G������k�K\�lK<Ǫ��r"�A���;��=�S=�.�M���c+0�n���Ka�AvS�G��m�TI����.@�C���䖦�f��k;O���k0'/*��'�K�0������;?�y�qlk�)���k�Mߧ�"��F�9��<jD34n��H�ˀ�*��Q"Z��t+�W�%��63���pѹ����H�K�VM�<C�t�o��Z�墺�
ɧ,�IZ�yET͚P�z ���O�E1/����7$�GVvT�n��F�&�L����@��j����ۢw�&)��pA������SQ1Q���j'EF�g�����o-�����EQ,V��"��vm'ME�F'���{=��w�o�~SZ���x>�+sn���3ܻPB�o,զ�/j�m�d!�t�m�j ����B"�R�<�.y�����>��V���~���̛��8ʬ�U/�AI��?i��x��o��5w�U� C��⻝C���o�qpWRNc:���v�ը>�`�XD�jh��W�V_��NH��b�1�Љd���&�&7D��+�Hݣ�� :Nc�����3&>�e [L��'���@	����K�R2�)�\���g^>U��U���Yr�|���|��ٚ1G�]C�n�D�'��F�@�� �i!�wX���i���)����r 9�F+�#T�h6X�P=��1;��uq>�9#�j�!��kud����;L8�s�&�! ����%�"�Y�B�2	��;��_�fVlu�tŷ�Ǫod�VTl6)��i,�l
Ig�6����k��@���;O�� i��V��-Z����Ih��vd� ��E ��X���-�<C���� !��n���2�߁vf��G���c[�$�3��n����Y�#�����E\{����A�ƴ�������)6��Y�%F���!P�5�K/�p9���l��IG����dc� >�����-��^��~{������r�}�N%��٣���k������w]��('f!%�;z�fCi��N�b�i�_��
�7�k��|/��W�Qn�6�W��;���&8�\�3,�%m��{�˼+D�奷���\����C74m��;���r�[,c-~���.�֓j���F ��t3��gng��-�cZ�uק@��cHjܢ���'}]����I��lV�����e�zNp*i��6�,�S�+*ixMn�!m���I��.��(���^��+��:�ax�[��wx~�_UOz��'�L��/���{@9l��X�<F�����h���/糛��;U<_ۉ���r��� ���5�V���K���3�H��ⲱ0�լ�P��m���{��!������Qjq�$�`�pM�J��/)V�p��2�wH'�����Zal�eA��)=�R1�}K%`�C����6�?�S����ߠ�~�Gb�J��t�c!����$V���n��L<�yxl��)�\���i�U��E[��ʚЪ�d���i���ހ5���N�K�c-�?:� ��KRW�pPU�)v~O@��������M�R<�Lk��t݉�F��nBLA�l��볽��]ܔ-�Np�Y������]Q�Rwᔟ���4M�3е��4a�B��u��Bny�-����/�\�byT�*����	�	�]�tC\Ѩ��a&��;�͸x	��%���w5�������5��W�8p.v���U��[/]旷�N�)������R�u�����t�ұ,o���KX�ͨ�S(�\"��c�n�㯩���ԡXr�tS����eޗ�Β�J��C`_-���%�}f�iRM烤��.{(�J5��	�d#�
�@�ݤʭ��N��Z�A�X	"��cMb�H��dcĽIdt���c���x��Й�|�L�n� �2���WJ�6�~m�#m��p;{c�ǧ��]�{I��y,)�=<� ��-22�i�(��ä=��ܰY����om��@q��ޞ�T]t+#K��v�[��]~�Ud���`�k.�����T�x]��hS��:{9�nA�K+�R>	�eEl�Nu��V�<R�0|"K��q��U?�\�Q5���zb��,��0a�ݭ��5z�#
!I6�����;��{L�k�a�Q25{��e�wH,R�H�D�h�[|	���=%L��jm�����A�'��ҕN}��"�V��a�>2 ��Ҫ��CB��z=�� j���ya�&kR�/ooKm�t0� @�7zDl��l��B�wHF�\L��O��l�Ko1�P�~}HN��}�"�.(Y��W�x5D`���EU��%o�F��f޴  ���y9�#7˫��d�:��g��t��(iZ�`fH^�X�������]K7=Y\��IE]�[��@�Q�@��ŝ&RYJ�6�\�I��X�/jjN�$W��ݺ�/¯17���d;x��D��@���9�t�����A����moF�7�7��b+I�߾^�Z��	hw�=�M�o�B���`�?��茶���h�rH�\p�[�o����ܼU���|�xQIͶ��_EM4t3�7��C3Dr�v�s�����<��n���I��� E�sU�\���3�@x�#�[�b=�-@�2W��-M@@����������})��^����d�ffeZ<��5[g��A�/חlO��<��_<�g�t�̹8�������䊨��\���H#{0)O��
��\lݖn���s�!�\�A���7��)�vj�C��^��\��Ms�f�lr����,��:�H�7a�o{��F �Q#ܟe�aͯ�"��]�?�|�z�>H��=�F�«��O���jR)��GH�����{D�/��Y��J�(���B	��"����^�&|u�Ҫ�	�] ��bi�q;*��|Q���|$�PD[G�E�Ւ��*�z�����͸06�E���q����l�uƎb-Vj��i̬��XX��V<17[�L��mh���9N���uj��5g�Q�J���q���@z�k�
65n4K6M�eҍ%���	G��E�򾫠:`����R9$�'�~u���_�>�>u��ܲ!9�ȩ6ьr�>�&��ۗw������[��\J�ŋ;�w4X�{��}��Y�U6'�L��CP5�#�=�3��$�0�>�O��/�ْN/�=�/I6�9��*��թ0"�kjsY��+��KY�C�AB�❴�73��wܳ���3b~�Q-H��
s<��C�����`�j�u��ؠ��V�^���
�$3�>0�l�/���y���&;��J�֨$CS˪;�� ��]~�d�2��	F0-�Ju����qjrF*�N���qu�]˔Y��)����b��
.��i�r�0���������&��9i_	�Ƀ�J$;9�w ���:�8�Ϝ�үo�u%
4���� @�.�_��+���-[ �6�P�9�,w�I$�C�ԉ�n�)`�"P��r?U�����%����Z��\�ڑ��Q7����<���q��n�hn�}��sF	��mئ��r��] r�xm����NF/�Z���,�ԗV�z�.�K��D_�^����}�T�=�4��er� ������ B�83��B���L�"�0����v�jW1c:�����II�������x�M���FQ��W�����ȱaK��'OE�l8햿N��v�&ŋ���{X�g �����^֨F��F>;����?���}�hK�����آ�yh,��#P�O�����"x��_�[-����(Z���F�t�x�c���He
E�͕�b8��u�ɭ�����*�YW�o�S�y.����N�ʸ9&�ˑP,�H�N�y�>Q��+�����}c��W D�|z��h��!jӨ�����	�-f]�B�X����V�l��]q3���U���^�޺�ٚ�km�f��l��Q'K����=�����Ugꍽqo���$I�e�W�\U�ݐmc�����7�<� ג�2�!x-���_6ate�$uHj�]?ۧ�í�A�A�Z�*��T ���:2@��N�B���,a*
�����a�U��]w�ԯ�iS[�p	���N�:��x)�Ukw��U!`�
��椭�7I87������<��p&!(ե�G���|#M�Э\A����G������z��/i�	��|& �
��/����p"к��^�'į�,Z^�kv�Q��y^uT�����WV�S;���3|w���
֨T��o�Qq�0���`8�_�0hW�����;w�u8f��R��־�����\�ͻ�B�r�e�1�qjer��� q�<�?���x��/>R�[xK��BZ��u,QYb�,Y+��o�0�T^	!d;ٓe��P^�}�i��$�c�0��jy��<���s�s���=�޹���d2uD�y��P�[fVU �/a�rh5#�L4�zE��#0�V�p��L�az���К��!_h���U"������3|��#���
��<��s�_��:��2�n��rʳK��3�Z�C�Ip���Ӓ!rZ�ּ�st��UՄ�w�ӝH�P�;&7���[����%�U�s�~<p�Y�aq
O
]���-��	�<�_�[��m��ßj�V
Q?��q��3>���,9�iL�I��~˸��b����^�Ѵ�����n��/wiZ�{�+<��Xf���j]:�x)�����p��|�Q�q��(��a���:r��i���#vh-0���Ǡ<�:V,�ʀ�#0_7&�����*�q�]�F��r�h�&�����T�����]�u�1�<���2��7�>�{�Ԣ�c&���	w��4�J����G
u&.��M��G����ڎ�6�صZ�EN5�Ϭ�%����)���տ׻��䶴$~�l�޾��m�ꋰ�-�Q*g�<�LX��>�<��m�y��޸���e��]k~~��28��@�m�X%gZ��lp2�x�^s�G��(�ҹ��@�`^
?�?l'�#t7�o��;
~s,c��F�ZWՎ�����3��fX�D�0���������2�fB"���|�5�M���F�����;�0���5u����jaч�����@�4�[r}��a��q��Uy.�R�vˤ�F��N�Bo1wϡ��3}ˌ��}}�ã�;����hR�HE�%��ʔEig&���0�[QͿ�;�W���؉WW�S篇���[yQ�a���}�t[�sY4n�NUU�������L�_/�o�Z�m�.�p�����Ғ�ө�1�,��"���%=w�������t�e�m��V�_�܁gV�)Y�nח���������q$<g'!Ɖ��l(�>U��i��Dm�ٲg*5i6��XLM���E~"�_�E�e��TMl���s5��I<�B�w+��c���<u����V�3�:���Ū������
o{ԕR,��q��-���3��}��8�ޮ�yʪ}��nHt�\�.������#�^�W%��-�n=9 8,&�M����YP���q{`>.�g�8�S��w�ߙ�q��2��򓿰Ar�:���fN�"a�L�Ӄ=#ˋ��D	�c
� "��A?-w���}!#�&#�m)�r�j�[\�)Ύ`�!�2���h;��;M"��-�K��}Y( �H�&���7Bύ��S�V�<'*Y�M�sJ0��F��~G/����^|ǧ���3�FE��ִG��V;k�3�i������C��+#�O�g��y�-��$��
�R������4��v�Nj�{@_ψ�uR��Q)J���>߇���r���K��k��b"Y��Wޟ]�, �j�^�F
�姖�z����殸ڄ���M.��j�`{LC�@L�N�D9>��M�j�M{pK6a'��m7�9�!���E�g5�*��.ÿ́dW����Ry�P��S����_����K�'0������}���<R�"�R�ղ�\�~(�@�c�ϐ�[�Z�Y0��X��`&nmWt�7�)Dy��Qz�0R�q=����:���EL�Q�С�Ɏ
�ӕ�j�*��{��y�ܼ\�e)ߴ���W�U���j5���3������`��\]'G_�G(S��BN�����_�PQl�,;��)���Nr��n�6����:mf�}�Q"+`ݪ����M)���(�nӃ��A9D�Y�%[Mx���鉿 �o4�z��x�1}ϕ���d�:K������v}󋚛�%�%��i�b��;��rЉ=xp���½S �����$�W�0��K�)�(��q�������{�47�V��_��UYc�^��Q��}���G\���e1�c��0�&fͤ�X�s��ۀ�j3��-7�"�(:U���S��U�8~�O}�_������2�mKd�<�D��T�mu�*������ot� _كoA��'��A�ӢsE��!�S���u��[}�X��¥Ԛcjuew0��3�ja���E/����C��c����s�~���{�;�%���k�!�^��<���!Sno��)x�e�,B[���ja���۲Նɪk*n���T�X����1lenͻ%�`&��.�
�VͩpEXv�͘5��/7�}�l�%�;{�q���!e�ir��#��3�i#>�#��(Sޛ҇��W�+�X2��"j��B�,�%AH+LUp�����;��(�������"TmY,��KC+^V;uul��Ի�n���w����Շ�����r_���C��\诫Sn�}��Z��Ǎ$7�?��y��g��!�{����vg�w�󋲎`H�@��t���c.s��������:�ё���K��*i�Mۙ{+h)��]��Ԫt��T��%��Z��6'�>�6�����;WQ��:/�*�~��+Bg@�i�kԊ�{�ڤvt^,쭃������ٽO/0�04˱/9���%H���
ѷ���jҧ=���$ݩ"q)��0����=q�#�(q��f�(��0B� 2/9��Z�@TYp,z~+�E�/8ܐC�(s���NE��:��ͬ:�`�N@4�v�p]��
Ԅ�%8��m���'�G�<�j����یa��#���h��W�� �z�x��3�S㽾��w�1!A�j����$��:���K�=�D����¹���3��,񉃕N:N�}��O
�d0�;.��Ka�B�C�"[R�o��B-J��'��o@�r,��o��s�7�Ô-Q�jt��/���c3�1��s#�j�{������ ��:�`Jl�r�A6�N1s}^W�o�*��䉣/�p)��@ruڃ��<T�?t��:��w�SO{�y��l��,�ʥ�j�L�}.J��k��/�������ڔ��b=8�{�� P��z�����c�X5������ݾx@��g)��KwԿ��ӷ'�"���θ
m������G������[�|��&�5Շ�c�<o�1������d�3�׼���;��ŉR/�_+i�y�3Q��V��솒�~������`0��UmZ^S�T-#f��9e�3zG�� [�A�ڷ�G���V���*lʆ�z&L�냶�v��t��ݫ�:�6>���6�D�:��d�xF4�C6>:v�"�1Z��j���@X|-�� %�~�7��H��&f��x���Z�K���(�]F]:�򌢺��w^�Z�;��%ݪXN��٪mT��-ۣ�h��.��
�r��1��:��I�Y�c�e5���v���$kb�}y�q�Ɖ1�v�L��r��p�|�s,on������0'uo"m���@���< O1��b}�(��b��Rg�Z鸡����S
���6B��q�Mȓ�<!O8A �DqJ�kyYW5v�3���ؚ��NQV��2;�(����>�ټ9�.yX0�]��cH�s?%NT��Ek�Q��`VH�چ,2No�/X6���j��>�,z�t�z}��.n��n�^�=����PJ������[��t���IP�@b�RA�R�r�6�ڍ>��{���>�����83NO����ʅ�7@T
�4*9[z_��Ul�Rɵ"�0e�{J�[󒜳fG�<��VZ�|ɱL����C��|�g�I�x�0�plt�>����}�K�Rp�"G�Ksw��3m���~~=9\vj^7����8\�z���	��5���=�CY��롵�G�<4�=G�.7bl�I(5��4��zK�.a���LD�\��K�F��_/�,��tuE�%�)4��Yĩ�����ߢߓ�!1	�ۿ׹�x����*����k�E����`h�Vq���OF3��u�]�Qec��>Q�����Y��߷U���3��#������C��R��im����u�s�YV?>0��p�>�,�
UVWap��=lk�Ya�^�������˨0��@x��¸�bd���35V)�Kv�Yg�یT[[�����}����᫘�4�l���[���8QKM+\�0y��fЮ.Kk��E�u����߆q����=��%tY���R�2W_�sw(p�ڸS.k���M�-q1
q��!g�]��ƫ�))%����nC/�[X>�������f��Ɯ�+ه����v�/ɔ���1�ٜE�Wo@2g@�y!>�F�J��9�ܒ�(�`��ݦ���������d��ۉ
��U�q<�p#v�}�Ǿl���{C+�n^�使g��!��aE�t��-YlbKπ��J��lz"GڦF��z{�&|@�W"���C/2p��a���(��#Mk�ōX��,�z�.�TT��3��X���Ԉ�}+4V�3�56A=��5���Z����QÙ���ܷf�IM5��c�f�6���T�k��!���zG�zb��xU+�{�=�✻D5ŉ�K�6��Ά�3�>7��K��m�-�T'���.��H\Gj��Ϗ^oØ��7&jj0�����D���4?��4��X����'x�ݲKr����5�bRZ����gX'�m32hӤ��e=�a�y3#�`��N�v2Þ_@�������H�%���x�2�s9~���:U�AF�x^����G�1����(<���&�O5ٌ����=2Pm
Mp��8`�����ec䀻ǟ2���)v�d���:�ׇ4h�1��X {���kI�����ɯz�t��
����<�%�����qf}�=�G���b����v��U!��g�9����Rcvd��R����V�]W�a���t�ap��xW���^ޖ���Rۉ��K�ځ�21x���&�~mcc��W.�bì{'�3��aϰ�飋�8<�/d�1��5��Z�V�`��$jg	Y0ה6�s����*ɟ�y�,��31��b��$��m����ǟ�bE�j��q-��Why۪�̖�e R�-a���2jPmɾ�z(�O���xp v�I��7�Ῑ��[�;g��Mm��Nr�<��Z�Hus_�H��uW�t��Q�(i�u�;	�ܽ,�b}8Y�D�k�Xmk	X�8+�X�b�*���*��GgM�"��Ŀ�@"-�u��L���GrckuI���侏�{IF�+Ǵ�5�1Qc��!�Б�	(O��� ���1Ο{�)�X�;�9�J"����w�zx���-r�n��?@��w��3~O�e��2�IE"�����+���t��zq��8�����X���~�����K�&��ʮ�C��<Gu9��}v��?���8Y�K�G����+���F5�}E6�'�R�qݪ����dЃ�W%�*Z�������Sg������|���?�X���c]Ϩ(m�m��˴��%]XFG�Ȳ/�r����������S
�XN#�����K�[�����I^Ώ�>�ȼ	�X���3T�N�����J�7�u�چ�u�"�l~������К �ǥ.�1G�o�u��=H��n`g^V��Ӑ���"na��Q���Ylٷo�Tį���VNz�i�۪U-���v/�_��fs�b��ɽ�h����ó����Jq��~��ki�;�l��7n8���ߗG�}f�}&}.��?�֨�9���6��	xB�I5��GlQ��+9^.O��j����5m$w.x��v�c��o��NЄ��r2�ﰪYF_~���^�X����A�������$�S��N��Z���o��}y� }��8���b��m��'*�q�Q�\"���)�vc��� ��ӑ'�'�p+��D���I+'�K2,�x�͘�!��	��|�\tM%���D�g6[J�V�ĎGl�����+Y|�ӓ�s9D� ���g�"���E��~��1tm�$��g�dw�m�ƪNtzEԧE����+��_�b0&��ei9�!��-v�)�D]z���X3�r��E�w`6�c��5�4!_�T���.����w�Y�����7���%�I��v�B-�÷?;�R_���	���ON8�1 (�B3l�������;�Z��F��2"w^3��ud�.�"��i�k��ꫪ�~��wY��!�y��������ޜ��M�9���R~��?�I7-�n�y�w��H˓g��[1	�?7��3��3��Q)������
��3��� �/���1���c��%4<F^�}��9��C����_!HS\��������;n�-m��hi�z�Afkğ(��R<��C��ɚY�ߓE��!����� ��R�����\�f�N�M��g�\!�8�O�q����ܫ��S�nL	i!���Y��P����٠��z��Lon��������)��1���1�c�H���|��o��H�v�Ԍ�~�)�\9��<�$�!�,��96n%8�������e� �Rz�Q#��.��l�kt�E\N�������?���Cey�{O@q��Ε&�����<q�����-����a��q��=�����LU {�ko��v����{�=9�ۗ��?�YRd�N-K�T����B:)x���p��o���E��"�%	fϟ���-�t���G�Q���Ѐ*�������S����*n��F���=��c�\��~��f�+��Ζ�Yl���>J����*8�:&8�6��ot������Y������o��V(pRA��m%��W�`HN��J2��@�KU='y��i��9��;I/�~y��w��z���XF��k�u5���_�K�����W_=��{G;>� v�@����9]�cC7q��`��0���x��Q��&*ܪ������jJ��{�[����*���8/�Bf��=���-��`�\I,��Y�I|�A����M�c����V�3�Ԁ���2V���jR���Ԑ����J	��G���)y 0:�߃��:�}#�=پ������qb��]�a�t��qC�\L����uK����iX��8��z��/�[`���YeҺ����Ƭ��%��Z�M��H佧�t[���[�#��v���y���%�Ij�r��u�/M���8������������p���l��[q�~�v�{@O}\'����ճ1.��o��^q9gPE�W� 7QO֤0�Q<ǬN������L� �\!>��٤Dѥ�F����5�
�_�rv��/�uk�p���J��=�{ �annȝ�<�ȳ���?~�Pq�s�4��U�Y_��ߔ���ڠ�t�[_Y=�?������	���4��`�oF�>Q�Ŋ�I��Q��Ʒ=�o�{Ή˱�����+r���滩"���%�?:O�O���G M������7-ң�x.I�/7���\�J3M*=�dN��u1��s\ j),��Z.���N��SJ�s�z�ۭ�4#jc�U�Q9����a�|dh��+<��w`�2���S�;�6��՗~Η;O�s�}#��v�ɑu��Y��āB�o�j�&�"-������9�P��`L���r���#)N�p?���W<�{�ͲD�*9�醁��6P�V�IY��vڶ*��ǡA�3 zv�7&vT�H�S�%�.jvO�{�y��P:ac��9/�e�M���p����#��g����ob� bȂ�[�٬#��S�;O�k�BkQh��*��s[ �I��.ɓ	(���*)�A�H7'Z�_� �k����0�a��p�ף�4ˊ����@$�*���7����� `i_���ɕo��4�1��4X̓���rjH��>��9K��s�`'����f~�� ��$���G����tN���w�a'/"Ia8��S����V�!�iO��n���:�,wk*.��el�	�� �7JHhի�ʬ������e#Cb�)~�3e^`����O��ä���%qI�)��[%���R� <��~@\���u�&��`f+ň65e+�D��-͊9���e[�5���b�Uc@^��4Ǽ׈�jc�Mv��;H�����͵�J��х�^3�V����Ϩ� �K㮕{����mt�0/{/�0~Q����JvY����}u��J��� �Z�p���«�ƻ
\�jM��u�@����������H)�pK��Y��l��~X��{���٩��n������@qEBe��2_#�Q贄��/����"`;	1��nޜ��[� ��[Xi���v���ѧ �C`�����������2A���e�*����і��ٶ�Py\1�
'H�ֶ�6���� X����P��qc�->]�Ȫ��T�Ũ���r ��<.(|�M��|�s���w7��fO���=���#�	v���~�!O�qZ3!M� 2�hR�����c�E	�V���%���$�TL���h�̤u��	"�
$&c�;�$�~R��d��)v⡢{�;�Z�@����������:K2����EE��W�P�B��b������=0�km�����S�.^P��fr)}�R�&H�ʤ�����~D.��q%J�^�5���^��щE���K6ɞpqȘy�T,�-������/��T�'O�_���xs����-����\��b.�5iƙ��b\\*
�m�h������v�d}+��vZ�e�#d��䢻��
�){��L��:�-b�l��߿����Lb�D�!z�l�R~"���{�������<��{�/Y�ɶ�hR��P�{w��A�H�Cr�n)`�RW�{�eRUYS~9q���aK�O�S@��1��.�ր��Y
�hz��9�;�C���#�F�� ^3|3d��!U��pY(_�;|��sqN�\������
t�)���F��]�_��I�X��4|����Ů���Cy�.�~%h�O�Y����7:�����k5}�(�.$��� ��8�iQQyAo���`)�M~����r�(s���{Cˬ�|P%�~_(U��*k�.�9�[<�<?���7�a��;1��b/z���?
Z�Ī��{�  �k����k�ju'����ٻ!�"�5S:;	R��[�-b����������_	'��S1���.\��%�;>�`c�+�`fg-PX�����G9{0P�E����͖�Ǝ���+$�>�_����G�pe-л���g�	��{�(9���tE�UbF�
Y�?tP�jo��C���E*oG�^��1C<)�@��0�� �W2%�����dj ������E�"=2�@WA�B� �7���.��GA�wTO|�:���Y�F�5b�3��#7�A�� �Kl�66�C���\�4Qt,�����ц��#��.0x=�u�4H�/-W��^�R�5ۢ��~�z��������&qw�s�(����?�s,�we>�=ê>֤n��P�C_��Zv��u�Y��۟���v�oVt��V�};}�Պ�	����I�=�<=��.&�`,x-��m�}Ԉ_�.��}�L~Q�2�(j�tD�+\����.���52N~��?Pm���׃�d��X���Wo[EAޮ%J*r�Ow&��sV<����f���a��PWR@,"T��vtŢ��z���G?�dU�q`ͅ��U���ҵ�I'G>�JȼF�N�n����d�W&����n�xD�K�C�O��qw?)*�BI^�ɍ]
�?�g�-@�`9�v�ۍ������:Kwn���W�A<9f�1w����>g��x��H�8{;U�}X�@���E�/>���o����V�k���DU�Ug"�%K�+�}]ED���U�~W���B�j-g�Ɒ��*B�t���3�"F��8���D����կ�|? u>��R[�֐��?iq��`*Ef�V��74�-����w�C��m�\�Ĝ(@�|�W�!;��="��p�G(�*��6��]�	�����~����W,��U��P�i�Y���|���������A�6�au"�DI<��\�3t1?�����}P�,���� l�2S�F\+�`��; \��ۀ��T�EѼ����ΩL}���I�z�7(<������D���r$FP��v�&yn+$�'�D�C����f����ީ&7����b�!7)tX�^�⪘�[�(��R��9_�\6ʩ6�%\��ץ�|�i�ƈc�$ζ(TL��Y?�O�s��;���XMkD�s4m�B{B���Kޞ�v�*�Юj���S�k����f1��Wu6wbx����;6�M�G"�T��6������l~	�=�t���D��6VӴ���Tά�_N�% �ݾVRb���N+r�t�I��u�da�wvy��|x}0.w�����=z[�!���a!{��? ����BeB�	���!�B�ƫ�Z�V#��j� ?�|�� �P��$Ue=��ό©ފ���N�<6'��qϯ:��,Yʒ��b���` �<i��
����p�D}���/E�� ^�f@�?�}A-��c�����z�9l���R�f�`Vc;9�E�G�k]��p���R�J��`@��.�쬑Ju��ȁm�9.�9I=z*Q�f5�W�z�5M�I.u�ZE ���M�Q;�.�k_����kQ���U�l1�H8;�;��#�)����#�@{���f���� �9Xz���.����֘��>��3�����e�K곁�1�s�8o�sY���7�r�E+�$��_��ӯ��ѧ������z3� ����ٲ��P//��R�����<u���H����7���e�v��|B�
�޲e|t�A��y��4�K��3�$��7(��;��n{ '4�_*�x8Pùo.�V�p�w7i@D��"t���,�BW�5g���.�w|����J�׍7D���R.`g7<`��]7�rF�B�ׁ�J�-��EV�U;��h-#u\����p/þ%��ZpH���y q)��e���qk}y�GO� �u]L��߱_\ء��Yd�<n�i����
lO�2&�b�)���A4������f��W��� �w�X!��4��rY��@n�1!�AW޶E�cE\�S\��e���A�N���Sk?�J*:�]��4��%vn��z�ŷ5W� �\�z�
sݗvC����t�L|�@ L�k��L��.��o��s)j�l�%:�46��zp+d嵼�Ţ�K(o�H�L�V�z&���[�Tǉ9
xѨ*���]�ʷhji�g��"����.@u�NYR��^lK��x�xlG�vVz1.no�cI�hE��v��\dYeY;������$���y��g�(�j���tU49g���*fg����q��gQ��C�s5�����}|ڴ�]�B��l�����x��ܕ�T��CeOY;`�̊��`����Hz�շ���\��ό�Ծ�� �!�.�H����?\<O�lM3bw�d]�<����Evw��74F$pj�w`� �M;��!l#��;E�k�U��>۾��R.������J�~���X�Z�U~~Z'��BwxN�iÝJ��l����V�)�ۯ�'2��'�q���\�{:��ZQ5[����s�M�^2$�k3]W���ɋ9���𼒵Ν�9Z�''�	*��K.�#ͻk8��,��t8���D���F�m�z���ƽ89މf�u	)�}/,*7 Ҭ.�6�:g}��w��S�ή{�А�x,���f����*�B��/�w���ZZR�v>�3�:*#T�u��;xK1�"�k��M�H�wZ�i����0�⤃FoP��p#3�
��|�L���:�l��%[�Ky%�냘��e��O�i귇�O�Dht�P�/~�3l��B.��RU.��~�řk�z��f֔Tu� w����<{����>��1z�g:ŋ�x[R�<4C����b`(8s:�H�;�@������ypG��5��X�6���k�1�|��k������m35�1|�e��˯Ky�ݍ6�`w��{td6o�'�}�fB�^R��Q,~�k��6�H)��l��?����v�A��*��g�s�b78���f��Љ*�m�Vժ'�����SZ��^S��WD�ƛ+WT�`��A@ ���6��u��w�M~л��a_�jpB�Y�� �ݏe��Z�0E^��7�@#کU�ϣ��ҿ_��*����_$'һ�r��}�~��M^P�C
^���P���"���J��\�^�૓e�+��B�f!�u�ޗ�eUt�M�7N�&�@�.�s�v�уD�{�[��ocB��#Î������c�2�q�ȃJ+d|]�����9�+wb����c��� ���M������Գ���sg�Qr,~}Sе/�g�+P�w�f�8���-�V��W\���~��J������n1�;2��\Y���T�+�t=�u5{iuX�����$s�%'��e2�q����۷*%��������}[2��M�Y�ڛ-�֓���0�w'�hR���,<��1ԋ ]2G7�<������F�������}֩w'	�����z���;i�qR.+���e~q�в͸c#�f@��Z�eq��f۱�+�������B
|ܠ�{�c�U��.\j�c���Ä��\��k6nQt�k#�ً?Fn�~��o���̘��^q�}��� �'��p�^�W+���4 ���h��͝!و
XNV(Z��蓟��~{'�'��ҷ,�v�"D�+Oغ��]��-t�D_R~�q�����Ph��N^r�_��-e�J�Uڢ��r�V�f����'�z#���7�@g_5��� XhKyHQϣB�9�Q~����i^�c�b=�J<>�p3�y��>����~ex�Eb|�+�_>���p����%@��?����~Qww9��\���3�� ��Vire틑���$ε�� ��3<��Ι�k��00�}�Y�]����[��4-\�
[��j���X��
1Vo�	�_�*�9F@���4�I��p���i�x���*5��g��Y�k��蝁o���5B�j�{�`�F����j���MjGE'WH�6+:��CO�F���`�&׊v�GU��@�������@��tiJ}�~o��IoIB^��Mp��f+�C>�3��ͨ!���J�h�m���K�cǑz����3��4s�����lE�Hu�f�md <�\A'�L��D����{w^M���g��-�P�֗	�ׁͣ��Ђ��ǂ���.5!~*Ë�'պ����q}�
 �7u�`E�M^�#:�n*��G��2�m��~R`5?ЫX�(�5��X�<����c�E�.���t1�&��,�d�`���k3��6�*����P��W=?�ƍ� KrZ�ؿ�����ؒ��I�r�q��»D���J�tM�b�<�j�mp0�~>�vXΫK��8aH�m�z$UN��~�{&um�2��Cr���1O��6pj����X"��o�ޯ,~R�;e� �l� ұ+���t�⢸�Y�EE��0es�qYVHw���L�n�KT*u���pԠ�:�&@�7&u!t���$��\[��Awm��_ܺ'�Py@ɸ����� �1��f���e]��_�(kR���n���FM����y`�~͛��}����|�F���޵��2��k�,�@>I�"��B�ǂk�#F�*)�bT�A{	��M�%�t���4�(��mG�-/��Jٗ}����D�wa���W�`�Uxb* �������*8w2ݟM�{����l^����$f�933����E�z��O�I��
j� ���5[6����+'���$�x�r�����qtzkmc�?�DuCf�&F^�sO�rk�s'O����oG�i_$��|��W��v=��遅�S3�FZ�9�d1!����0�U^(�"�UA�H>eS�H���<�tQL�|$KeZ#�T��e}M��J������i�I�x�C�cQ������P��!O��J2;�VSF�ٱ��ݜ��"q�[����� ��7~���4�نϷ}�O]���)
a�q�f�{6�Q<���y�����g��S�FnI����$4�	B�[nA���Ěl?�&�2S/J$�8�]�v��v��V���p �\T1���ў�4*:�vu2����0 F� ��Tp,��[S��`6o����buG�ؔ���$(Q�+l�*���M��Tu̶�G���'���k��*�0i�`%�F��#�D�x�0�gia�噐�֗+[�1��ئ���+�4�r�%ǥ*��	���_ȫ7&�5P��J��A1*~���I3e5�D�g�����lUߊ��dWζ����$������+��7��/m����r�e�����sy�m��]/�70�69e��t�O�9c��B�R�����jچ��mZ�P�/�o���Km+O�4Z���|*&c5�w�Z(��Uږ���<~�r��fN�p���`0����U�{��v�i���c������>���_!OZ{�(
I�Z]cQ���5���-v�:�����g�W���
�a�U�{�Nw�{^��e��aMsJ�s����ӊu���c�~\s�yJ�g���&����K�2�&�zEH5):RǷH��K^�>�P�����~B}\���D� �� �����7�N��}_�oo}��$��V�+JJ���z7i;��I��j��-"x~�|-���HgbnvT-ǲ��(dK{�F��o?{)@QL��\�]�]9H��'mz�+sk8�j�%qE��Ee`���K�RڔF�5g��(mu퇹F��i�-���v�o�yq��-AF�r�3s�E��9ɪek��g�SY�,s[#�*�����l4ٺ_�$N�4�c)K��f�CF�/��"��
�6�4�W��+��(<:����u�&��I]�Ď��0k�}$=���/����C-�4�7��k�P���`8��8"E���)�@�qY/c��>�{A,?���f���4"dǼ�o�������l��G�������?`F��^�Zyum�O4ױf�'�,����~�wCUG�n�Z�K��K�~��+�YhQx���D�8#|Z����cLK�����o�K����j�]6Z�F�S�G��V�c֝Ȥ�WQ�'24Q��rKԷ$Mθ���╗�C�jS؋âق����v���cv�~+�0�}v�gE;��t9g=��is����<�)����2`�fy\����|nU<��_H��	:�\H Z(Y�$a}�!�c�0�Q-E����W�$�:��`AE�+q
�|���:*�{sb��Zxf�Rr��/\d�
���7E)��1�@���.T�Wa#3qp��&8�������E�&�%P�b}i�5����rη�N�	����h��3��>j�^�\��wB܅�S=���W$n=��1;�r�w�v���M=��e�:���Ҳ}u�Tq�_�F�_Sj��dٽ�Y �?J�'��=�1D�}��{f�z��"�������k�f��s�ר魵1�j�j�� ��P59��m�D:�3�@���q8N�w�� WA�?@��	�'0=~���މ�|ڭ)���
��v=�@Y̖����Nn�ƱꐑZ?#P\��	�jj@�'*�ݑ6�غnW���Z-D��	$�������]��݋�Cr#�T�{؃�߮�yX�y/�a~���A����)ٸ��3#����-�a'԰,�)���1�K�n��r��4Ɋ�N��@�'n���b�E�aU�������5�"&R3�H�z�yᩎ�V�soO��<��8��>W���$�q�pn�룔�����"&0J%�˱Y�����>�Qq�r�.3������nD��`��$+M�7#���"3�B�xV���HbǞU������|��_�yա>�c�@h�����_Y}�ݻ�A�]_���H���Uh*`wN��:z���롃<��}\�f|���ve������C�7&����_����EU��xCС�J�Lm���+���`�/�
��2����k6[��;�v��.���{�#��֪�h��K�Jճ�[l��u���[�2/|�9�^��/��9]�W�+@變 &&���o�ĖU�h�Cј�5����l���1j��W��A*o�'�w��T���")&]O ��bm����[_H"����b����lq�ܕ�J��@�Ow3p/l`�!'��aW�����XX����x'h������?�Y$�X��ɫ����v��%�y�z�Ԕ���D�a�e=��4wW���O�e<�]/�h�|���2ooƿiZ:>�m���pN�+c��-/V�	6
^���͵l#jA ���$�z�8")�+�i�r1Z-����
�cB�&a�6��fu�߼<ԴUO����]�KO�4';�&�,��\r��'J!*_����Ư>�ne���MV!�D�*�XH2�vo�V����a������M-G��:��.>�lH��z��o�[�X��=���c��ܧ��M��]P9_p5?m9&<�(�jv�J�҈P<���㳝oqk[/�nLte���|�k���i��f�jI��6�X�Ja�gw������͐ �ӏ+A��U��<V�Pg�XLupO~'Dc9\�k{X�2m����(Oyq�,��6�7Dbk��험 �b��~�$v�Q�)�S��+��PA$�	��Y ����&�Α�oOl��7d�_̩�f�;�I���G;n�}G�ˏk#���W��A¸���:�A�c,�`�����;! ��F��G�}}��h���A��î�Q�\�B�i���Ogf����vn���렟�t�����M��e}���F�k�}�8����ҝ�]�iAZ�{t#���������������b��8��y}o�v��wg�tj%�{�_���O��3._i�L�[���Q&��[Gz�be�MX�/3y�P�s��e����;%��7�@��fIs�,���>_h)�:ʃcĐS����>�Y��l��c��nlJ��D��� ��UYIw�̂�����L�C$�v- �ȳ��"�2e#3��4%�IwQq�� 3yX��Z��D�$g����p��.������n1o�z]ht����n����/�7&cN����Y��%q��2��9���r׶B�	e�9@��E8�(O�+��0���K����m��#�m�����l������S�X�z���q/�
�:�4�j���H|����I�Ϲǖ��̭7��E�hTr,�PZ�I�@�͆�2�q�G`��߮�[f�������:�f)(?�������P��t4]d��p0Xv�ѣ�Y�Ө]�9of,i�٣1��ʾF�/0t�^J��w+�m�1�ʬ���,����Ԫ�Ȳ��=ʕu}.�ؼ��>ڐ�t`�"%����X��X�Y+����$2,�2�`O�thN���-Y�,o-���_�	8����l3]���*��CQ�%L��H::����ͥ}Y�Շ����	|'�����kq��C�pW��s�����eJ���o�@0"	�g�cɫ����._L҃3���}��,,,�����v���R�g�\���=�zL��5ɲIΥ���gW˒�VR<S�g�Օ{��o�s.�b��<M)F���e$̭�c�hЫC	��u1�<N�0�G��!�M����N>�i8i0[ϨG��j),^9)L֙����^`���Ե
'ݏ�F�C9��mKf�i����B�/�[�;f��_�hC3c2�.��tC��ǝ�4�3������0�\[�ˍ�/O}��e�����;�.��Z^�v�u����4��G�AY��n�7-l��=c�n�T�Dc6�w�Xߋ�~���@���m��@��$r�|��>*�Q�2u��ҳ���(�9�#�?��-g�I�z�C�2b�C�~91��-��k��n]{�x������{9lT�Ջ�ϐ���r���Hð6QS��g'�����ٺ�>��U/�$�;�J�!�ɘ��}󄞫�{9��w���p�<7��-���a��!��R���Jd��I�a����<e� �AK��!�R�y��k��e��#�Ͼ��sT��u�p�	�=�iz�:�#�s̸k��&)R9�^}c�J������;XyX��;��Wa�#͸U�V�u+z��G����| �3�j$_B��Ջ�@�:,v��X��Q/��@��Eފ��L��)Ί^��RF3�U�����Og����lg�'R��j�A�mj*×y��S�d���@�:�^=�'�ٷ1V�⒕a���E�����ҍ��;.[���������7'խ]��;N�ۚ�<*F�p~�}YHd���u�@:--g��;���������扆�i��Z)��#;��{?����>�%��4����<L ?�di�ޭ�	؁ڌԧ	�����U�Q�^}~6�'���{ڜ��	|����y�d��A�f�6+�\O&n���ܾ�:��p�}[=ֽy��b-�&9�Q�0ǅ�>+^g�6��\�yy	S�XB�����nN~S/*���D���O����ox���q� ��^�*��Oٽ=Is�M�>��4����.]x��]��YRY��I*=M��G������z�\�e&K?u���
�/^[W�n����b�k}군�*���R�c���NI��&o����C�וY��к8���a�� ^ן�C�$��c��`ħ��$�ٚ����.1L�v ��c��^���:�����lh��m����̛�^��Jǅ8) *��ᒅ����^�|�]�{!�v;·��Ƙ�?��g�����%'h���v�A��� ��	}9L�hu�@#�ƿ٤���>��f�\����w6�n�F_!���	�Sܸ'��<TǮ���Dߣ�׉�rp�қ����^���ޡڴӌ�#>����u�I�D��~������S֎����N6����jl !يB��e�-��{��럃v�I�C$*�����
�m}T��Q�ә~����MEsɔ�;zn������٤Aw�âe�ңu�1r�C'������}�XƇ~�yvGx'��w~�%�Ҵ��8�V�;�|��CGq�c�x��2���/��`�׋��{i�p9��Źn��W�t����N,�k�#�}�R�=i�o�R��p�7��̖��k����m�-��5q��ҭO ��;���{s�ýF|(���洭N-�����l�_���!��
���e�W����N�`�v��X6���G24�6]3�R%UP�
�3�O|k�*4wWP�H��C��4`7��$����OX71	���z��.I����uw媵��W�	�����"L5sn���H:>HNZ;��.Y[��:s��NJw����v��f"����߯ŵ��������׫�>���� 4�~[��;Deo���>�Ʒ$tAHȢ�E�[���W]r�� ݀.���Js9mfˬ#��
)f��HoD�57Hgz�� ���o��D��g��z�*�H ������6|	�x��
=�U�K���olQNq��Yϥe���b����̄���7����Q�'-IE�f��_���Q�Ѽ����ϛ���Q��ዞ�wS�~�{���Պ�u=�=R�<�چ��og�B�@_g�"Ӧ:�u.*dg?ŝ<d[s�d V�E��J8nx�4�,aoڿ�z;�Ǥ!<J�'��A۽�0��n���
��$5�Ook��1��&Һ��<O(Z���Yt�i}�5H���t����-OV^�w\|ymF�a�e��4&�F�~�v���| iV�8*�Le�*�v�5<X�V���-`b�͓u�����Kp��E�l�v/��CQ�ٮ��L���L�}|smB90IS:�x��$�ɑo�y$lwU���^��&j�q�$|ȃ�f�N{�L�uJ��ޱ(�3ˀe�$�ck�&ˑ�ٖδqh^�"d$|��4,Lm�#��b�wJ������p+~�.
>~���d�?�Ŵպ���A�S	��#4�r\�3�ZNA�|=q;��&��h��{�]{C��i\|���ݐ}%�αx
���n���lC�0֊��e�س�����T���H�,��
1�Y����e�c�گ#��u,_W�67����'��@����+����-��%^��eF?�*C@��ɪF�3��*T�.��φ٦v3�[�?p�[њ�Æ����^��2gDG�.��c$X,�ƅ��:5�k仇޹l��{�%�3���i�>8�$�����Dv��B���VJPh�'�S(���*xJPϖ�k��I����h��|�OV�"��L2ۊv�*�M{�4��7A`W���5��k@H`>}486�D���M�	�GIJm��~"k�u6����a���ay��?)�����
2�pg~��>�?p���,v�-$��2>y�MBA����R`z�P�q�h^�/.����<)������|^qxr�y����drR��i���f(�~/x�V?%��=�W*��:VL��@����N�d8A���L#��χr)�pyvM`��o.�rf�0�������Ҕ f�����H���$��+�"T=��.,�Zd���k)�%J�Ǖ
�B�(�ӪPO-�\n̏����CRs8�_ɟ��2�?n7�&�Y�Vm-��ϣ2V��(h��P�
s�<�����}{��%o��(�%��'V��Se���d��@�����8���*U(	�c%�^z�ya��2�^Y> �j�u�jѧ�$����ruF�5�������<Z"U��,[~���o0�1ʪl<�?�e>��8�m�NO+��R<~�d^�I���~�����^=��Sȯ�� �s�]oSU��Տ�q^�m��(!� 8sNN�e���ܜB���ܳ���S
��c-a'wF	���+���<0��ZE*O�z,���8�-�0u���f3C�*;x_��'�8��WQ�z�����U�i7oqv�[��,�է�{L�ܡ���DrH�#?&���Ա����D�u�!�,3�r̳�"!�SkF$�g��"E�DV0je���]T�_ĐX�
~�ڢxd��6U���HIg�O����G*5O*'	-���gl�Eth ^�K�����
�g���8 �˖�5|�"]��9�p��X�[�H���L�n�-[�:�+�ӷ�^�_rC��F5� ���^��G7�W,8�63��MBY5�7S�<�Q�A*��TO(Գ%by����粭v�'�a+���>ߏ}�}����ɳ
N#A�O�Y��'g��#!m�%
ܑ���`�TB� f���^�4�W�_�O���2���ZIe�2�[?�����'�(�DX�!��G�k�8;wda������]u[�_Zb����̤D�:��X(�Q�kcQhS�~����3���O0��pwDXٲ�[ ���{b�G	�6�3 9b�e�#�������ݯeM�ۼM�K �O���x�D@��J�B���J@��dm��C�X����Yƌ�O��~�ڽ��+�u���0 '�1�U���{s�SA�����n��;���>?�L0�%������Is�$t�˾Ok�� �ڮ�*$Z'�?���ݮ���.����l��P�T�͓\�Y������W,�Pc.w8���*Ux~��ڱ��dd�Rd8�_�=��P�-#����WP��H��G�ث�y���L6�!��de��|8���9���G�����:^w)�\�?,L���kV� ���PQ>�c���>d�	eu���}[ZB=͛�]}��֭
��M�	"�<mXB �����O�f u{���
��6�[衮U�7�n��/d����	��*�8����Y�)nw��)ۀ�ٝϵ�>+��~��߰v�a�|ʞ���������"����|�ha�S���?\���}��~�<zٗd��{s>�U^�E��3�s ����,{�#_\8��dk]go܄��a����3#���e�a�<�����}�d��Ϭt�	�P����0�W��.�qe*��.�J��Z�ˆ�枣�i���	�����M}3�@����B�48���{S�vl�.�
Kov��-�':��蜁����"�8���zv+h�6-4@�߰����1:_ŀ�
�nqü�f �}V:�q���]r��:�쁒P Ժ��Y3?�]@��ӵA>5�mm����]+��W��!����|��W�n�ܔ7����#PK:6Q��/B^��kz����S	,3�f����T��l���i��="[��-��4�:L&�rb;��$ᜢE\V�n�'��/�0�!�r	��ob�zÓ����g}���/��Q�Q�RcovWG����a����@�Up[=Zê��
��u�A�i��6�X�C��x{?i�$�D�s���,u���6�huZ�
9�����5Ϗ	ӑ�E|��چ1~g�st�ˆ���!����a/���������L�/���.	R�E��*ݒ^Rd=Ѽ~�ghma����,91t;��\�>N~�n�YA���&il�,n�v���R��ϿnT�w�Y<�/�������?6��5��S�d���"��1���4�I�8�S�E-�p�SyT���H�Z��W���(��ۙ,��7כ�֙��.��:N��kC��C�p�'2M�T"�}ԁ�"e5�]�;&�MiB��.o��I9饽�,���&m;�g]G�t{C8����[w}$^�k���侰z�(�������X�`�C��`��j�ʏ ��O��VJ6�@s���M6i�3�5��"z�=���9�e�Z�P���r���P��]�+׊>z���c=P쏛��c�})u�������C&5R�ڼV�PQ�N�����3ԉ����6����G2(�l&�s���������[�l���w��2�[��H+؄�A�U��]���;+vU��)bGy�����ޜ���:���� ��4�ä>�u?ڞ����-���:����ޫ�k{퉺W	W����{�.�ϓQ�U�>�D�à�Qq�j����g��nx_��ci�ݙ�I?���`���pF� �������犓U�19U�Zӽ�uJz����[H�u���3���N�88���!&�ůr�p���d Xz��!m�j�p�]���r�|~sSwvX3�x���
n�tJ�跖��x�t�82�=zE|�%(�@�O��d����WoR}�K�݀�������A-ϔ���$R��9T�z�B�rG�0_j'�pa"�倉�7ȹD�@XO��.K�5�����~�pTAj�'�_�s�~��A�}Y� mh_�/Ɍ6 �=h�b%	Ɇk���E��q'�il�}T"Y�p{�k��t����;m�>M�z�'�-�Z&�f?u';<�M+���<1�q�����
��4���q�m���i��WK����B
�l�ԑe1�w(@jZ���9���ξ9�\2���\�FN?��
܊������?��`�A	�i��ځ����,���Uu�Oy��ql����)Y4�wK����=��^E:�1�>P����x8?ZX5�^���4��W8�U��4�ډ���H�$?�&���S�����9`�ON��=�p�݊ ��ޭ��`�����콩��������Z<��&2�g7_
^7�ߕ�>��"�^t`�x/e?��t�q���� �x".*y�C{�Z퍪KpB�Ex�C0��F��3|pz��R�=T$��uvZ�U�������} w�ҟ�����0�u��a��~��<��]�A�9��{���Yk���V����A��*#���%lʤ���B���6�]�!�:-�X �̇t�&P������~��#T�r��$x;�D��	��5������n'￿�&��V���$D��	CMp����b�`����^Ӣva2w�]P%�S�wQ�|A�&A^h�V-�M^ ��B������?���qLҕoV�������)�c�*��������D�g��n��l�0I�0�$�����E���tA��7o�n's��j7Og��A�Uo�&I�Z&�o�Ӕ��%� �e>q^����wr�m��c��/k#ݨ�5Je��٣�'|-A���
��60��` ��|�b�H''�9�|T���n��σ�/xCV�%�({�����\���-Ҫ�T5DՇ��ն�'�f�������=��a�L��?��RU-P�*r��n�+4�zQ:�M���x�>�>�����D�aI�ߗ���N�O��㾆��?�7�:-�9�::�L\��p�7�ֺ����X�u?b����p��O/;y$gkW=Y�K���#���"G[x0~,
�<����S}y ʬ��Ϥ��+_w��8f��2�L��AKj�9��<�B|v`�P�n���.y%pCT5�O<NS}��@�|!ǘf�z��G��G-:��la�?Z���r:�9z���!��4F�벬=u7˴���gemOX�8ǧ��בM�=�z�Z���=Aϣ%{�J֮�Q?43��Z�eF�`���mE��D�R9���[�p�6�q�b9�7��ma[��o�ǚ�׈q�ű(�]1���C�8.��/�u�d�
0��S�����͗����x��x�Z�����<um��w�����Ȭ�-�C3=Mi��cW�Wp�8�CF�Ҝ��[��φ:�����_\dTV��?-;}��{@�������0%㝦hɲ�[2 ��#��6��=�C���X4���^N1�pc=]���>
�C�����{�6�k�8�vI�5O,�1S�B�~��0�#�5�F�Fg]M���R�{�h�8K��H���ГӶW�c�7ڷ�����߮��2��3�D���l���3ƌ�bn��ܟv���aܽ�����a����`�z��dE�x����U
ɽ����1��u^��mo���"��܏��-���9C�ij��(��-�"�K=�ҽ���y�R5N_(vvi�*��j¯uA�k��h[{_�g���J�w�g���>B>'���N:��`�*�zR�D��4m�[w��¦߬����<\�eެ��rst����?"�������1��o�_�K�DT�4��a}h�`H�O��6���Nf��u �%�ߕܵ(����f�	���J��L�q�nzq?Bu����uڻT�6~���{D8�#۽�&��%^&��p�VX��<8��0IcN�Cc��B7��Kk������2�lr� C'ym.k�(S�B�%����E�Ԗ��l��h��R٤��ș��p�u�]�n��<��<j�ҊU�N{�^-�5T���Ź*�P���w�]G�������z�7�5;�~��sia{Q'_U��~q\y1����K�-��2���D�o�p�?������n]-����W1��@RX�wS��1ɀ�T��x�f\D8��.s�&$߬ )��ȓ��.k�aK֩�hё{n����h��bN���oMr܇���,�,�XNCT�p_�k}����Uɬʡ�k�̊��L"�ח�>�i�4f�����l����<[���e��w)�+|��s6#/Uq���V:������%���83~f%,[Q��R<��ې�&	9��T�Ƣ�%] L9�秌VMU�.P���>��,�Ζ��d�WC5G�7�Zţ
mli�waM"E�m��8˹8���'yf7g��6ZP Gxt�z?�ְ��y�2O��kko�io��4 f�}S�V81A��^�����:��4���yP�|�HA4^�����'n����7H[�E���O�Qju�Qg�r��齱;^��z��˞ɷXj"z|zq|w�I�V��z��CB~�節�;+I��96�b��J#����q�F&��eY�q��h���}�'4g�2����礣<7H㫳~UI�+~�*��m�쎗iq{h��)��Gn
��]"�!����Ԧy�o<��ӕ�ۣO4\&3_�
�VE����*�����>2ߢ����.����0Re�@�y��F��ۑ❭��ܣ�s��\��76Hk����¨j�P�6,s�h1�3{(\�n6�v^�k��}��A杓|"�"��]�AI�	���l͗^ͼP���M��C���p"-]�D����F�)%��8B6��!�%��]Ϝ��8����E�;���j�m�2MI�/���{��,��B�Ƙ�&��)�(�^ΚK^^Y��_�#,us{|�]4�|��)U<� �Kj~%��IF��4�t [��2��VE���(��Yv��~�|��u�I-ipr��ԧ�w6�Y#�[qbfjyr�����в�+*�#*QǢߺn�\t!ץ��u��/��W`!�l�n?�ʬ�GÁ�����k����ZuA�ʳ��@Ȟ�k��K�\F�ڐ�|d{�Ⱦ��3|P�2Z��YqP=#SZ��Gg�{�����_��҄JB+����=�n8靧V�5�v��Lu9󖿑���� ���!���gWw�l��abPS*����k����_2�6���Tg��Ɛ��q��̱�J�ş�Uݓ�{�h��Mx7��4΋{i�fFz�ǚ�1lh�S3��Y��e�A���=U�E-��Y�����
Sj��;��0�cCǷ��kD��<UB���{{W�\���Z��;�I��r}P�grʊV���8�k��6N���wי���\��׋��wf�����\~dK�]�5V����|�_�G:NW��B{��?��6��d��ڊ�.�槚�Q�������v�䈪�s���B�O ��gz�'���*=}կ�!���m��8?;D�7<��>�']!�����U?5.OQR`��>�_L�>3�R����
.�o񘑘�=B�WE/�x�:���v���7^�<�M�����@�u�-B:��K����A^��ff���, mx~��ۿ�x��������C������
�o�# �e����K
؂�%c_�Y1�+3w�	��B�&go�J�gLo�6)�`gC������a'b���x�E{�?]5��3�Y�QRp�����J������a0r�����xPpyg��dsy�.G�^�?�F˅��S�?� ��|ZN����z���U4�p���F���'����o[)�����p� �l��j�;�+���P	�q��+p����߇I(Ar��%0��YH�mQÌ��T��ΨㆸΨ�o����;���Q�� ����r2 `�r�c�����q����P�K�s�I����V�ݘ�|��;o�kh��K�9��x��񰯦���s�_现���n�C�DO���B���ԟ�^S!O�n�N̰ho�O��6�I����h�\f�;,Gw����B���>�.���2_6��UHӬ��.ֹ���Omi�����̾`z�ed�8)��]�l;s��Q���3 �.(�����]z�:��@ݝ�������
�q"���[Z���fo,����/��.E.z�=ˁw�7��S�7���-����j�����DQ��1���iIkW�L�4�P�sp�5˩��"/��Uv����o��\�99��,�������i��FK�Wx#�9�AGVV.(W/�+7ڻ��l%T�	�(��NBL�C��xЋ�j��yL\�p[Uj��.F!��?��jʢi�^�#��*�$� v����'ۛYN�VF���~����4Btx/v��J��������r'�d3�طb���e�dK%��Cw��Y��2�<LNY��b3�4��֒U���S�*��g�-,�Fi@#��l��%����JԷ�_��Uգ���)�d�wr*�5�5I.*�p-ӓ��Ǭ��Σ	��R�]�I]?���MW�ؗ�,�ɬc
C7c�����&�	X���l�u��k��6��|<{�^��d"RItf�-�X;i����'��'6���G{xꊲ��p����"�[�����N,�� �]���O��
��q�z~�ÜN'o�/5ԩ���Ǘ��P�%�{��/���X�b�T><�/�~��=s �5�c!�B�O�L��f�aS������`+x���vf�<��[98������GW���6Nm$�.�-<�Pe�V485�W�o��(�<?=w�|�h߱��œ,�c?����|2;fｋ!��)F�A�N����	u�O�j��A����'Qi��i1�ߦ�%�v���A��"?�	`�JOx��ҏbQ���g���2�"�u�f'�m*���2�)k���6f�H�/܉@����ԛ�ܻ�ʌ
K޺���S?~b��n��f���;4�H��o%/��*���k�QT��/u���v3���p����r]�a9�1�cB�]���zu��	ޫIF�©#2�(���R���r�)Ԗͷ��:��}��cy���Y�)q(+��+��Y���[dȴ%�,Z�~���u���[���R4
D�xy�+�|���?��f��Ĥ���/Q4�i�=z|�7��*/���.���ug��Z6��CЃUM�xݟ��oA_R�u������M�� 2�mW�z�,
��k��5�1��?�����J�n���ڂ�W{�k�ž��}/�n�']Ԣ9���۵�l�p�*����#C!_�qoiw���TpB0�)�ٹѫ$�s>�#7e�}�ڷ�f���$��������W8l70��e)�ß~|��1��N�����$G�ܽ���+Tk!3�!~����'{��"n�,!�W���h�<���ސ,��M�@o���0���:�j��&7! �$R�ke�ͽ�@���!�H��r�ݿ���h�-_��-�j�)pվ�*F֊p�F�`u�v�$?��m[��~ٜE�RB;N�D#�F�@�;���i[�Jӽ��5��oG��ĞykV�L�����|A|�}�7��fb<�o��vG
Gڨ}E�0uY��C�88��jCHO3���ſg�a���}[�����n����۲�SɎ16g[���$˅�;c�y��0��Y��X�GDkA�\Y4�Z�Y����B�W;���*��Q'*�F�w��=�ϔͯ�5�O�p�4lF%�b�e~���T�H����8c�䎲R��܉����^3�����^vk>������;;�x����+iOa�f.|t�H����S��ytˇn��E	�����M����Ux>H|(�O�P&w�0xW7��Aȯ%���akm%��:��ʻ�0��7���5ot��(ܥ�����R��Z�/5�̄�^��A{R�F���d���t�$h�i������ݜ���p��k�56�n����~��Z:ߋr�%�S�m��ClO�w����N()h�#7p�V�4Dk���/�Q��C� )��_��ـ�����b�\�E���l 鏙dDA�E��J�<�*�5���C��;
�"��2��¢Oq�K�{��3{�X�y�.P���������~L��*�E%��Pi�o?����h8��u)~�b6z����,M��]�Ÿy��흙�H�7 vEV��6��uE9��y�.��=�9"A+�}R�<P���ď�sSqy�����X*=K�������ɺmP�:���o��s���s��0_RIf������^�d'�}I�8M��Ne9L�T�k-"�;Aɲ:��d��W�|8j`P�S%Σ�	�qK����/��bv�A��
�J➣�d򑿍�)��*fU E�&��Jn,:��-Ol����=
��mgx5���ě�4iȲ�JC��?6�wΚ�c��k+�D_�g�t�����n�&�-o
ͻ+�����w�2d�0�aà�c�Oܮ���F�U�o_���?C�����:�Ӝ[�;)P!�W`���u���� �I�`u4_�ڰ�t�l�ȯ��6��<�R� B3�h����!����U� �x�?1��qȭ;:�Tн�IV��Ԝ����['�����tU��?���becs�0_���{��Wf8��'o�LB�7W���?T�)�is��'��v����xB��شxu�-��]��S��Β�W�`�b{w��	��Wx���^p�4�4��$��2b�ܱt�l7S%� ��+B���N٥���ȡc/�A)�Ydc�,��"����q�ç"���&��X��M��̚��a�m�;IWK�ixO��&-��8�ϊ�DD���P���m:`�3��ғ�t��@[7\4�a���B��O"=N="�D��Em��r���F�m�ڱ���+�R�t���4�ԓ
�@�N�ܮ'�=y�������?D���hv����w���*^��l��BQ��ְ����s��F��%�x�eX�R�lڇB5L���g��n�jF2���:�2LFKyJ����7m1n��
w�k�D�8�DȾ�5|�z屹����?#���]8��(�#U�9/���K�R��bY(n�����Ter�9Q&Xn����pk�lk����bHd�C�}8��c�mrvk�l�0dL�&���ʗ�:��i��?�{m2�G�F/F���z?��gƱ��-l��ݥ����~{?��7U��D��W��꼮6���)�$��&�)�����Vq�.����3.�K�k�̩%$R����J���x ?Ie��\������~l��$%�&�R'��l�9[�L�6&�� ҃�Q��{bl��X��X&�i���#k2��e";2	xzl�8����֩j4U�@��(Z�����4tnA�M���[u,�ŋ}���9�^G$Jː�kϪ����{�� �:�6�����qvś���7!�c��{���[!�G��}�	�O�������n�_TA?� ��w���?�?%%�ރN��M��2��	t�i���	����f�vX�����W0x#y�O�u:T3�ۙP�
U��\_����l$���#���x���i��ka��iQ�p�&������O�'v��I�Wn��"5�|ӿ���tȫ���M����o��U@?��jݷJו��[]�H�P�U$`.�m�lB�#��f�be2�}���z^ ;������&��\*�][�ъ�ֽ�zi��Oֺ+27�N��C���A�W����c��Zbd"�ȭ����n~"S��[R̽o�!8�b�\�� �	��j��P�~E9v��54)�ciy�a�*+���+N�k�˓sߝ+>��K�����l��t^K�h\{7���/-Yl�G��0Q�����D&zj�.I&�|Ȍ��&_s��ݞ��4 ޴��
_h��,�����}V(r�ڔ[�>`��蔆���A>zk���0n�_(�ْ�m�Q�q{���Eof��g�t�Ը����oe̓�>��UAC^�27�҂Ŧ�oȰ�h�|�{f[�H�=yx�j[[TkY�=�-�X˗�IR��ѫ�Y�[T]#<�"��>��H������W�� ���\{j���kΈ-��c1 �SX����+\��FE̜�ǻ�~=���t
L/�w�gaW�v�Ce4��A�S����W�������3=e���ˇ����y���Q�8�W��/��P���'��c Q�lQ�o�D���ψ`x��_�!�@jWC�W�y���Aщ�g�<#Ҹ�t"VW7Z�	�΁��蠖�����2Z���H��H�Cw��Mo��f�n^R]A����v�����.��F@��fU�~ٚ�,��V���`��������rV�ԑ  �{�'��i�\���W�!-<���0�O��v*�����g1�kIɆ ��� 4UȖ��u�~�5fL��y��i�2��p��{J��פ���������hH��0�2c��[el]�b�x.Ư_N~>-pP��ƕ����[N�Y���"��-�*�VC�O:b�^'E6�7���9�J��*�z������`;��5v�Mgj�����lk�2<-%����i�Or�������Wg�M�r�����"�B����H���i �Nh�����!V���	㴆8̐���⌤�־�G59�JK�3���;�4�2jc���YÐr��2���R��n�����R%���E�Ǒ9�X���aYd��b�?�`A��^��0[�ǈ�a�6.I���eGѫ�M���5��W"�&�Y7�ήl��K��A�]���E2��2d�Y����3ZI#oPE�F`���#x�%�Խ!���E��4�V/�Tfބ�G�a��٥���m�p�S�h)�Im#Cz�2�C�*�"�M}A!����;�Q��o�8��޶0�(��+��>�l�Oئ4h��ʻ�� [)i\[:'���m�l�u�xQ�����#bqBS&qq�پ�W�u}��
/_\A.��_մ!M�bn|��f�����u���~���ĲT�I�������7��Q�}�v)3*K�&�5�ކ|��;���X)��k�-����3���m0�d,�uW٫0�)���!��hF���c͋����v"�>��P�v�GN��dq�6� �5xCr�7T�,k�HD�b����3������I�^k�����DztA��.���C��^>��V����:�(&�f��o��q��{��A���g�a�/M9K���|�"Y�#"���`�� �����Ozy�GZ�޿=!�����)|�X�1��2<
�_۪�EV�<s�������i#�� R����t�|��0o���s�0#�=�b
�{��E�s��6f�aa�9��l�-���:U�1��,jZ�à��������뚍7d1?������^f�'��_�G�C�_}�.{�Н�_M#I�8����]q�ՓYI8�r	(�č#Bn�*Eq�s�Zhn&���њE��-��t˕�D���e���vv�Nyh�?U������Sd���[;cΉν�zI�>~;I��M֛f����V?�'��Ui��7=�&��V��3d�N���]W�?��� Fǎ����Ѱ��Owc
���0�_j�?]%��b��2�ц��(-+�Mb���m���m������zH��ӓ�X6t�~rA���*���5�����LLĥ�_��}E#S���Q�l���`��8bS�H;`�j�[A<e�ZsP��8�W� <M�s�-�^�r�7;?�k,�A�pp����.F��R&��H[Ӭ�vk:n�Ʉ�}1��G�v=D�*�]��)G�Kn���(&>7��o�2A����'����CpXn~V�q{Wf#HX	ޡ����K.6+	�P�X��Jeބ�K�a.PZ�$�܂/ki��AIa��&�ݣ�!��4�[\M���%�;'�����3��4���C�dpw���·�����]u�=��W��Æ�#��A�>sq~�5��o�+��j�xkL�cA�a词�4��A�Y����:�3l(2E��@���{"J�#Ah�i�:0�S?��H���� L!Y��:�F�U|��pG���Va�eJQ�'7��7�������7Z��S�e)�_Ң����f��Y/,�Dѻ�I�V�=~�%TɸV	�������3����R���C�[��"$�ٌ6�v�X�@��ݟ�ek�##�gZ��.���q�5������ ���*���_�)�>Yǐ��C�.�#m��n��!"�9���ə�fA�������e�#�Kz�K��N S�0�XD�U�#���Q߆�UT>}�m��*��t��q3ej��K^d��IM>��Z�b�z|�h{��:"칡�u?�p�x�G&���}�k�G�{�v�!eE`
dJLȎ1�g�RT̀Z�,��)3�3*h�Ei��u=�=�M�~o�;̮�V̇�X��-�P=n�"j�d���n�G�i*�σ��;W
eeU�������Tg��K���YF#~����Cb�ŷ�@�!�FC��o��d�?\'M��ۉ�;N�!r�&!���&�<Z�v���B}�#
�9��@�H��\��ձ@�S��WRD���<���]�����K쓾�X��KԌ���3��k��n:���S1��O?�����s���3����F���5&QU�=���l�O�(Ȏe,Fm�ҡT�c����^�c��i(��6P��`<�P:�����( cĴ4�*�ʓ�灨X\��̑�{�Ҳ�'W��$&����:Fk������D"���Tۼ�w�Hr��Y���Sf����
d����}sbB+HT���*8ʩ����{�Z���U� ���wŗ���I]�p]��+������d�4������XQd~��:@�K˩m��?�8�%j3����þ���uB�V����g�}���37m��'�4{hD��/���ξ��'%GF]�������O����G�hH�v[���G������ea�b���tCR���:�N���)��_�L@S�H��y��Ǐ+>�P޻�(_0������w�u����娴���q�1��Y��@�3�²�A�V�C�7/�X=��c?���D�.T~wF�$K�Z�w#���x��t=���`�G�h�k�#�i������ 6w:\N����w�)!X�^��
p�	�M���I��eڎ��{��p9IMg���֬A��@c���k�=[h|޾^�4��8�Y�#q�9.��
�%��!�1�V��������M���b�ߛ
n����U�Uydw�u�� ��ʷ��t���;ΉJ�m"�M6��i�G�����FW>�w~�c����ϰ얊���<���is�h�P�Ǥ��9�ٽ�����E�� L�4.�en
�ԧ�7�������
d��>)p\x�k�6�B�=u-�Y:�-�Ur���yW���̬>oϥ�BV���*DE��zy��B�
�Di]��U �`���%o�Fg�L���kL)%Li�����������2�����>E��A�bT&�Z��KA��%�Bwd�r_e<%j$ƀ+����ί�h>�=ّH?g�o���Yˍ�_��[����x�!���e��R?��h�E{9��.�P��jY̥��.��-���n�r�I栊R���Pk(9F�w|��-@h��Gb����|8�{=��Ю#�b���ڼc�#%]��))�� ��Qp,�K��m^<au������[�C�_G�����jr��zm5�����l������X�f�ey�>F�GRMj$�n|�q�H�B�m^����S����ju^��`$2j�[U��Y�~���v�����zB$�"|$+���� "�{���FCA���#��l�����,܎��X�l�6%�y�7��3\lܩ�~�)���G+�-�x�;���g^
�A�-�h!�F��[��0'��/��覽��,���Q/�T�w����ug��<X�󎼲Fe����]Mtd"AE��>8l���[��-�+)�h�]S[r� &T\��u�,��L�Iw'�ʲ���#f����O�P5ٮ�2G���3���C�,2��j���J�����n c^4�o�ї��d��e� �|KIֽp}e�gX�K�L�״N<D�
;�h0�zc��l�H��2��QpԾ�0��|g��}oN-��+\���}?�qQ������(cBBU�?6���n��8m>y�}��&�������C%�.o�Za�Q,��o\��-�e��Ә*���t.��͡RJ6���DEjL�KS��+���5s��.V�'��P��_���|[���<>�F�?��.�	������[��g��t�%�z�>vK#�8��}>l+�2>�	J��S�kP���F�G�kˍى�\؄�	m�;&{l1���o���^M
78_6g�Z���z~ �;����֥����f���kF�O�FZ	G�!H�m�@&�)����cN��Z"�4�^��05�q�����2b�����翲/�`����޸/P���ǻ?b��̚��:6/����N���^Q9�S�Ch_�<v��ID�t����w�x��JK��)N+�9 Yr���B��o;!DHb	�����r�=F̂c�,ʆ�T��7�%^HpphM<�����Cm@D��8���.�?4�q��ff/�m��ib��Sc�'ڒ|�
��Qew���xj /o[�/�A�>����S��m��R��.�xx�a�#Z!Nn�!�N�58���6�lU%����C0��-���X���%I84.�LY�v\ޞnѩ�;X� ��.��h�
���u�B�ڦ�;���<b7RM:���Ȭ�+o���t�`Yr�U��3y=�{�������S�!v6�N<��_X�����j��,l2D����X�5#�Ȭrz�w}#x@�;'�k���#�7�/>������G�����\3�n�fy���b��.�i)� ߐ[� O��/��ꚗy����e5�uU��Y�Z�Z�.��U)�@4e�eA���LT���!�[���<��v�	f���B֨�`R���F�;�D+b��f�nD������Ğl>oV�������L�&�/�����v��86׭&AL�b� �asdb�L,uɲ�4�z��8*GH/���f.���n�T>��DN:��$���uV�V��W�$K@�� ��<d^G׈6��3�x&(�X:a9��ܒ�t�������Z����*Pޝ������n�;u!x��9~�d/s]���O���E�5�c[�{��A엔O��h��V���ׄ[�l�Qܕ�id
ޥ/l�H���2~��f�H�<g�b�< -
�!h�rO(0.�+cP�(\�ź�w�i���[�����6/J{H{�dk�4�j�܋ۯ�<j���X�<��������k�D��%
�1s�p�L:��YN-!7s�+�o�hiÁ�J+ ��<d�)����ްI6�q�Η	�����?�lg�d��Z�Y�7�E~̝n�߸��kXm}e1�i��K�'�m��|�n�N0���ݮ��\O�帖�Hn�~��\�A_�&�+��N�����!h\��%���Gg�T�l��jx�7=�e��a���@�jdI��j�pD+��Q(�%	E��#u춣 �
�H�H�Cn&����TM8�H���c��-?@�e�{mٍ=��p»Z�Ɣe�B�Mb}!�����c-�>��%؞	:y.�l�u�U��}�a�Z;H��c:�&/�*��;�S�/!���`�NAifb�,,6]�"hq/p���� �L�A��Xÿd���}ƕ,A�%n7C�*$������I�<���͡eTޭ�Z!�t#���y:�ƞ�y���FZ8;~�q�h#�:�\�FE����<���:5Z%�RIO��܁%�sWK��.��]]ś\��Y���\k���z�:,�U#�N{��!E5	�.14� a���p�Yi���|I��lx�m��6�� R�����]�`'3+��侷�����y�����UN�`[)K�Arnl��,I6��d�mq����KN�☠�����y�3>m϶N�;J�7�	b1��pv�|K#t/��4|�`��#���}RG�94j�boO��LM]@`�Hrw�{��%?�����J����!��K��uJ���[���*iL�7�3�/�F�8�-Y�_sP��Y���KӴb�3a���=�<;��Q&r����䩳�5d�&�����#j��c��8	�72��˭�=��]^?�ݎGԳ�;%ѽ��bh���8u��E��!��}Ys
�8_�3ٓ���h��#F��N�+���"�'�6���h�K��k3����(�8��T�)&�y7J
�Ilx�ԶR�5Gu1��e���~ɭ��$
}�÷(�)2f�`Y�٫E��#4�}C�u�K�KD�Ma�O���ְ,�<�K�:Y�l�m�$�6"��0#�N�"�'I@�j���U26hZ��'�}CSt�1�1�nR�;��3��/����J��/ى|�[�?q�$Կ�2�U����i�J�3D����r��r޻̶�>i$�0%����j;6�$���I���K�����ތ��G>~�;�o� ���M�
��qw��m껼�L�X}g�e�p����6(Z��U��BGS(�,��8��R{�L{Y�?�|9�ҧY7��U�X�4ɠ�$�f���p&���o��!g��Lͼ�_7I�b`<7�C��~�N;��t^�7�4I(���\�T��\!�4���G&�K�&�#,k	v\��s����FNm��8QƧp/��+�A� �1���ƹ�~wa�v�2"���`���6z��c�6<�*O� �[��p��i���Za��.��Гߘ������� 	a-����]-�gh�7�]V�7Q���/��u����ysO8�\��-���n�$oeBe%�B5ͤ�zXLe־�s�M2�	�x8�^������v�{l&v�X9Rs��L���r�f#�Uv��ʸ����ߚ׭��h�3���u���<{\ᘩ�	W>����]��X\�
A<�-�Xam���*9a�*�C_o@#��6Ω-����(��I��	�a�9�����w�����=-`竨'݋;fS��oak}/�'{@>�'|u/����ɑ:���9,X���5�^rrp���K�~��%�#���-���7�E��7{Z�uH�Uj�=����f��X�05=����]}�>�P�{�D�7K��E�pQIW�F�Ϋ�zh�d�'���Ϯ|��&�����v�$/$2�f��ܼՁטq:L�9o�]�c(�1�E�gI��J�e�DB��#����\���)c��2���I2^��Y�-�=���O����g���ҞK�U&��箄�������bBO���^}��y5�M��eQ+4V�IO���^�/>oKc���%N[ˣ>�|�\���.�im�-�sNݬhy������`�K"-A���Z�2����_~^�E�w˽  "UbTb���c�E�]��z�S����H�A=��LSO��{�,˥;�#\Lk�D�z��=EE���"��x���6J�[�=���Pό�X ]n�3)�'���74�q����&RXp����=�G��AFK;�k;�8G#��w�^O�Y�-!�i;�G�4Y���⤉[�?w }i��T%Y7�]�RY�	yǾ�M��X:R6>��e�Ug���W���m��Ze�!mԙ�&@�o��*;�JC_����x��ն(�wƲ~d�I!�� 4�[SO�J؂�8}F)�}
(f vq����|Wi�����e�umEbИ���\z�iȸ�9�m4�V3�0���R32�^E��הK�����5�p'}��A#�
�R�zD��Ŵ�b`X����
��)Qi�#���q˅F9(:��<�ERLXQ9c{=%���@�#���S��!��g���>~�+%�mB�.1%=�������M�X6�"X?��4ظ}�Y8H#���g��Vr��u��ॅ��H��8iS�Z!�`}K|��������)Kww���!Ο��)bu��93�	��^�=28��f����
g�,�7� oI���ة��8%;���R:������� ���g��G�7?�^�L�,gG�֏\��T�հv�=uN"ZB�������".�*O>'�c�9�8�z��g�jN� 3	ALdZ�om�K���zNr�Z�i�Y��|�w+��T�����&�+��V�(�OJ3���am��1���)K�o�Z����[}Zz�z�������gw���@m�_�
%�K[+��q�s�� ��:��|K�$�'�9Wx�4�������Ӊ[ܴɠsU��T��v���516"SƯ��(�C��B�x���t�R�T��o��cB�N�۠���)�7�J4���h�K��&����J�TvR�(<��v�5�᭢e9N��%�tX���e�G�}�����u���?�c>�������sn��
��1�^��6_ށ�ǈ�@�%�l(�c�p�bk�7��/emx���[M �=�����#���ȲcZ����.��İ��3�v���W��r0k��C�J�����n�:��_�"�>>���+Ү1P���P�{���
�^�5���ܘ�����e��*��}X�N��<����{����+�y��h�x���+K�O]t�.���E��w��[	:9\n�����)a�����[�#4/���j�kh�c��b�1+�s/�6Ú���߭,3�~��χ����9
;��F���)��Q�u �A?Ty���T�c��w˭��b��D��vX�3�|X!�[2�t��'����d�@�3��%�QD�uM��V�e�h�7π���j	�1�Êm��_ � ?����F3R�O����3W@�Ep9��Ca%w�{�p8a_5	�Ѝ�e
?�v�W�,!Y(���_�'V�Qd2\${�d.K�q~��yQ4/�]���Zs�4���[���3t�}�Lu
Y.�m|�_<Ny�p�&���9���s�Ȟ�;H?S���HB��_��l��� ujz�ƾeT�6^��ܷ�	橿wdg���^9����6�M�f"�EիJ�q'��}vaY��P���X��)�M���Q�["ݡ��e�F{}����F"���ȴ���:		�(�cZz=I)�d t��X��?�ʼQL��D?�ylQ�fQ�{\G�)��c~�:: �	�K��V;�ȏ���\	����ѧ~>��E��5ߋ2�>��𢲻�p��V��:������3�~�����f��#L1h�&��Ȭ�����?Xh�5�xt�]%0�tIP9�մy��o[�mV!j��ȟ�U)�M�g�f T����X:�����-F+�G�m�ͧK[��6B�~D����x�|����;��0N��t���湱��Ǝ��=(NVnz܆�����y;�����a	�|>�1̸���,�)u���TU0���ɏ���N�����]О2�su��-�G����v}X�{�Kޢ��w7'��p��]>l��\��C�4��p�z�V��h!�.Y�ǝȣ����[쏅��cXK�7�P���H�}]fA���d>M�'�΃��֤C��8l��&�Ӫ[%��>#zx��u��8���h� .~��8|���1:=)�+�����9}�C��]�v�JW÷�KY0l���>��A�AX\�����{�d���}���Q�r���?���T*����(��A���K]��*Zr�yW���/xza�S��H���VM�o�����U�Z՜%�8�9O2�Q�����U!xy�D$����suNk\6��IJs�����Q��lK�G�b"�_���B��YiU �=��S�䮼��=Zʻ�"a���oA� )B]�a�.�
_u���_ڊ
����X���ۺg���{c=H?M�/a
ML����G����p��݇U�R$4�3�,S5�*B���'��)����
�/�pd|j�4�A�#8�.|X�2��O�Ʊ�K�NK�_�_s�o������&"���U+�.��|�Ge5v��w���w@��7�K+=�$��̕���
Gp�	!`�E���ǥ5م8��fD,-8,G��DC@m��D�/L?�Lع+T�#��U�1���d���6������{k'�~&"�6�=vC��ٹL��"vq�9۟rׄ��&�|�),h�e�2L�6LW��gU�dǶ%�4J5�2Q��(:N�c)�f�W���|���'�O�&ߦ]bJ�=1&�Pۤ�h�����g��h݆k&�G�/vb�ڜvEi���(o���)�9;ݻ��AM��OE�E�.|�%u��� �ҥ852��ж×bh�����A�����%*7�T}�K��]4��?+��X��}���D���Z�B����c�g���M�R�s����	w�pr����ݴhֹ�?��j�]��o����w� ��L�o��蘑e���/9L�5��V� ݝP2���F�	X���M�����<p�Α��V��d�6KJ&��*�ڲ�`��eqW( n3k�q��,�}�{�O�L}H����ׇ�<~�R��1,+�R�;&f���h^��ߚ�m�M��ڎ]�p`����j�oo���z ߹�G���F�:li1)�v}��/���8����	K�B�������bɘ9���{��6Po�I�jh^��إ(O��g���`}���J�T�b-m�xS/�p*:J�s���_񫦂jqZq㊻���QzKv� ����t����+�kO�"�D����^@������e1%���s���ݶ.C��>�0V�o��?�8rȢVC��Ա���94�6�n�n�[�y�,�S��A/B�����֨2[�Ɓ�$#P�����,K��V_FB�B� G�G�j5K[9��\	X�X���Ŗ�^�P���p����
J�*9�榿�\s-
n����r7� �͠�����t��!�÷l�}u{��"��G��*�F2X}�}��s�g�E��_�"ujh�W�V4f��<Wg䥶���.������a�Ŷ�ñ(��]�0o�1<]�n��b�ɛ4�7���+ �T{4Dh�3�m��h>���;��Sc�H��~�`��%#-��Z����������Z$b������ͮ�L�$�/� <�^<�[ۙ ��/V�W�Zvw�w/��׵T����a:�2�G�P�1}��V���yb���~��?�t��[.yO���g�y=�"��4��Pަi�S=%��(���V/�~�%��/Cv*��#p�6��p�k�����M��޼�㤫#�,��\��	bozx��`�ո��o"�C�I�ߛ��TM����5��j?�D"z����z�ơHN� 6ҕM�Ɣ=Q���~ra	3�֦�N����W&���6Y���̓\����[���4�Dߗ �!*s�a)�s�cD�d�s���ո�� �@�5*ʃ>�{ƕ�B�ڥT��q�oѵd6pf�*���s��N_Ew��eB�f��~YԨ�B���}uu@x�`��zq�A�U�����I��,��������&�|�V��5Ą�e���F�����G������ի��Qgt����[2�C�m���ݖ%��
���a�M�6_��d)�'Ä3焵��O����[�od��-�\R�(S�}�����kS2���	�p�8:�[w�[��\I�c��r�I��>�e��eT4�g(�]*��݁�A�*���7~�&��M]"=1��"m�ط��5�V2Pa{O�6��V`W�q2xӀYI���i=�L��eג��sژϷ�qj`ͯ�a�3���æӜ�FW4]�E�+��,@�b0Z��"��knԈEՕU(o���m�_&�K��M�ki�����X�[�6e��ӕ�]�{�|9,Ȣ�s��gw�b�O#s�Η!��+�6�V��4������]�$\����DIX�~�o�:(D�:�e���J��Z��q�i�|:�a�>�!�fK�4���*�<���0�-L@P 5�ҝw;R~z�U���e����`��[l�)8.�$� �r����ԋ����<��^�e�n�u���O٤b�&�oɣ�d	K>C钙a�r��F��}F����Jm�����^A�� �yCk�
��U*h^v�G��_3#��)%⧌@lT$l�ߍ�t �&d�ک�G�:`i��A��c�o8_�;i��OQfq����Dl�g�L�Y������#�\��m����5d�t��]ǮSm��|:&�'?��U|�$��3��L�^���환�B�K�b�	�8�g0�N\���Z�t�S�BB�h���̞��1�M���p{�Q�	�"��s���Y��Cz;Q��2|��EP�gB��FW�a�&B	�Ȁ�bd�ˁyS�<�pvp�K�h5�ź������,�����cr�?�G��%_���Vo���+�380����A:Ș�V��;��*�\�E���s`��[6��}|��T��&b���`��A Bx5������c�E�o�m4�i���$��⑚����%��ᐠ���l����������'R���Дs����b� �I���f!.У��"�%����SBi���A���Y[5�Yv��O����u{R��q�߹P�&]�$�W�?%�?W�%�m�*�B����c'%q��tMqw��?���$����K��B��< �1p���J�1��xb�-5�ĤͰN& ������G�k�.q���ye�a:%�Ʋk���$�mMe��u���Ũ{�|(�����xŬ�]�b(Ŧ]�Y�	F�	7��#�P��Ԭ*��l�vSS����s'?�&��>��Bs���1����r�;�X��{�b�>�J�pr��r%g/~�ڬeE����>5�mb��T;��Z�E�}��CC8�ٴK�/!�����9$	�J�x��bg�5lo�>Ծ?b����~�͖5��+��Q[��Vi���q�:h�ȉ%}�T���kk�Bo�_o	�ΰ|�4��8A�_ �W�����{�?Q���܌Q���A���N�C)b�$�ո��p�_Q��ƞ��[��x��ڳ?+nx���f|�q�_?��Z��v�rܥC����j*b����v���m�9f<��.�;0�xǨ_|~!N������+�ŏpN����X�k|�WJ?�h뭏U�O��|���d�|�%JF�k�3�n�/�ޤr�N�6��v�s y�-�
&`Ż�s\K�C�+ͺՃ̝�[�!��d{�zS�V�¿H��\}tF{�˘Y���Z�!U�_��{ʵ^�r|�ԏdNS���ٛM���߅�d��e��j�/�?%�D0I렽|�Y�t�%Tr���}��j��OE��be��Q��;��A�&s�@�z#�^0��Q�R;O�%�N!�l���ӒV�HM��HԿ�ژh��^�K<��.���+�[e�W;-�a:�d
`��0.:O�E���&~��]�U�,;���.|�.;xxe�-Y��/v7���M�9���q��Q�D`�,� W�ul�e� v���O��3Ƒ��|8���e�Җ7�:v��|n�t��SsPw}��|-��/_e��~��|�����sܜtg��4��M���6h���WB�?2x�}�Vu�Ӌ<�׽C���� _	�<�O_��[!�4���yK4 ڸ�z�:Z�e	�H0��~[XK�9ZS(�	�4�F�U�%K&jڴf��`&�ɷ�۔��$<S;s��4��Q� (��Ds�0�o�l?2Q��j�U����tK�5\������=\�m(�[��ه�\�����tB?Kyg�
F�~��~�s����"�kYT���U��՞Rs+�;5�6�*���F��!{i�� ��Y�S�N�����������E	�Xp�����-?���\!}b� ����DŪ�=׵W�����尤�����׮�G7�4ʖ7�!'���yE� ,�}��&�܅k�?��J����4:��܏�e /���U�<�12!T�	�6���*t;�#��].6k����Y���fw�M���b�z�f�[������6;W�,��t��ޜR�,7�&�!Ƈi1�Ȉ�O��|*�рio*1� ��U��W�w���+Y����C�W�x�g�T�:���[R>��SU=�Ъ�=zR�8��ɃhK�a,蔱�*Χ9�[;���c�ø�_`�l��Fn=�;��+D�M�]x���@�3���0-G� ��4�P܂�e̷��L�I�A�N[	!l��؛�!���"q�OB��a<A-�_�8���p��ˁ>e"�q�N�MX1ᔜwy��iq����	5��	�,�$_�2���1	eܑ����ex�����W����F!�Yw�5y���Te�L3�k�>E�����~���m\6�q"�х�`���㤓�.���U!]Y�ɫ����w�8lm-֝G�lDƃ�0;��f6��O�����3���T笽ETW~��
˞��C77v�1"� ߗ��A�"���S݃u$P�5��3b�����Q�g+��������@��Y�2�d��#�:S,-�HnA�
F!,޻��R+%�f�~�;ڣ���]��KK}�K��~�U!,�B���r,�Z��hr�7�V#�u��6he��F��[Ea�{�U�����`耜GِVٚ��hu�Ɗy"��H��-��}�X���%��+R?�wd2˩N�����s/���U���Xw�q�Rlh��4��k��a�E
�����ZE�MȜ쨸,�ܟ�b��׳6J�0���2�NAL�!���`t��!�)I����b�Vm%�} Q�'�-�n�Rp���][��Cl	ɳ�
��:>S7�����`�5t�I�G��{�n�(�uH�]��wPr�̡�bB%���\�Pm�"O2��OR)�i��,��"`Kk�&�4	S��K�X���n|�>c�����Di�T�ժ�Ż���	cXѮ���h�1'$�������\���m��^����?:�+�#j毡�qeQ��L+5<Q8 !��p�_�*5a_�E���x�������-3��p�f���j���aBxk��ëi̬�s ,+C��21co�������Yh_�������t���]�`�����f����/�3�z�ĩ<�%X�)��F ��قh�i���PՕ�S�P+ ����֮2/��W��M��P�>S[�iĝ̣��=F?6^zd�-�8Z�8T�W�vN:�"of\���phl�:�a���}91M���"?�73o]�mT��_��o�І��c�(����%s�32�����!`�7+�� �I�M���?��t��؊~��b꽔��Q�F�~�eTH�ж���S������)
��)�ojJ����[Dr��w��	�k�m��!�3A�Di�O��.��WDd���+�B��2�
Z�C	[l�eP�VORk�l=���6q�۸S�X'QMBL]������^��7#S����r~Y��!j\eq*vY,��GOoy�}�V�7��5v���E1p�� U���+�3�Ϳ@5�;L�}�z�'b��+���_{�`���>	D�ɞl\��+W���"���C+nT�_�>����Wr�4AAF�$�W4G�ej���{��(:�K�)��^>��}���j��о�1j?7����I��ۉ��E�� Gkן�H��X�m}/8(�5�0�B�߂�B��Ԫ�R#�>(-U��&�7���X���K��_4��-t<s�iB��\o�À�Z"�2�I�K�%���J��U�����ky ��=��Gҕ�ԝk=�|�ӛ���`����"���eJC�t�%X���\ӯ�Un�(��n�.u{�ઐ�wS.f���;@�9��~n:����UR���d��f�M0Z��^?�FX��j�x���d>c�Kw5��Y�tEk?~�j�g�+aǧF��ju��k�W��p �pL9�ŉ3�Ƃ�f�MW߻Fa�'��T�/χ\/����.6d��K����C���������'�p�=�'5u���sB�"*�Zx"t��l���$>�xzA�o�'A�s=�G/�;P���eɰC�B,%�0��8�+��LQԊ�98l��\�l���5+ ��i����e�+�	�7�x��IE�f�
6�!ċ弹Z���P�����M�78�=���h=g�����7�-��~���	bBm����iܱ�jE��>ׄ��i+cMf]WH�tG-e��W^1�fnze\ �?vp��iO����**��"(� ��@n�;hWV�Z�յRx�f��/,���7�aּ��ok�_��2�Q�+Z��jYŰ �h#F�(���0���C�`g"2��ސ���XV�ro��Y���M�,$���{Q�{N&�7���N������'e|�@CP9�T`����%��5�>j����Rw޹��5�c��Ts��Ί��͌'�_M�H �#�Vɠ4'�j�z����2N��S] �t`��I$,�؊AI����_�xVGw�������	N�;y�<�yU-�D�zy�#����=?`0 }�t���?����)2|J��:%1̪���V�Ӟ@�e��WC�������3W=y��	<�ɯ&�JϜS���S���ha^���_�D���ل����45���Di�Q����/2�}+6a�0�f����~��6l�H8#�wε9�+�T���~�y�h�s�a�ܰ9u��:�����rG	3JM�]ռ[,�D+r�}+v5_���>����q���3�Z:):+���~�K��\ȃ?��_�Q;O��'�:�F�]�J�#���m�7@x�"ET\a�P�,*�L�-}������]81�<V�����d��a0[6K���?���m�n�>}�0���N�I�-�I��Mo~�O��S�l�2~O�Mtt��|aH���d���n��������>��O_�d��Jm	s6.�����M�z3��5�d1����1E=?_�V=Z�g��4�e/��1�� &����Z�U��Dz>����@�����|�3MӬug�OƬ_��� `����h�PB�s+.�Q�R;��?`4_�@�')	����S[ȵ��ja$ G���5����YH�	r`�۩��#���ŗ<$��#b�{���B|e@��i��u�U]�j�R�C����}ejp@��j��i�p?t�q'FXF�~��y��8(C���v�{���b��7�z��ۄ/EB\��.��[�c�򀜫%Yy��	��ԝ�x�2�)%�S^�@��̎QN��a�e��r�aݭ^J�͇���<�s��^=�t���A3�'#m��4:xg�u��q�.}��d|TY+�r�Q�6Ƅ{.5lg�I��
���_q��m]��]ؕ1���¶&�(�zm�%n�h��ؗ>r��p��l5�6�Z�B��k�	����2]�#�ݨ�*����*�����ŉ	�'ԢY�������8���z�R7�Z����iJ�	�Ma[y�g�����ך�����e�ԢvŨ������dsZ飝~��Ί�*�e(��o{�.��6f6N���[�!A�z��Z��M��1?dm��S�6�O�~��Qt��ZO�R.GBU9<�c	�nC�m�*�睟�~ӳ�/�=l�um5|�}��<E`�n^�T��a�y*0cUg ��죲��r+͸�,��Hɖ�l� �������P�=;�l���Mxo�Yٓ��egN3����O��>�g���ء��ﺰݳQ�OK��$y��(CE�nmR=#]2#^��[!݂�o��<����JȈ�LzV��5�c��s�� z�k��m�x~=/��x�-8��e�4��v�a��k>���|�a��*�"�����J*�O ��(�R/@\������������!����D1d�O+%���䶯ψt)ٖY��I�u�vvڔ��q�mW~�lLA����P�\�
�O���i�p�X��t���P����yD���i$]�g͔7�2;H��y8r�S�v��@	M���G?��Y�Z����8̗m�4������Q�Q�����"�v9���F�M^�;c����
 �	�qZ�'rr߰Y�9����M#Ja�~+}��Fm��ܿ�m[z>�zi�*���&;>HS�e��L�U`)L�k����L�ߚ:��3]7c�G�[�q%���ʨ^F��<s�8}8g,/;�� A;�z�X�'����#[4��B�C����'����aT�=:��k�#j�a��׭�����7�_KtuX�Ϡ���T7���W�q�� ����-V,����(	�*�F��t���w�f�� 8_Z� 7��4�-�x�ַ��}��f{�1���+�0n��f�q�^��)��B]���J#���A/�v��O�Ӊ�n;�	�IYkO��&<�f�q�I�p��y���s��T8T����%]����;�����UD�>�%����$���n�C�SP�NA��A�;�k���~o��?�r�yf��9����h8�`���U�Fg:��U�)'�_?���B��E��$�����nQ�Č�V��Et:�fa��{j��k�2���u��S@v~|�9���vZz��9<s̪I�������u%󃥐��CʩԎ�=&�@�[󠊂7�O}�� ��
�\z���hU�̝a�Tb1�)��}�4�Zl��$��Ky!��vq/,��Y>Hv�9�)ZπzX�C���B�M��u���c�@(�M�)���s-9m��q�V�H~׾�7��(��k`���Ic͇���`�T���kM�beP�@M�yH�V�&~.�����q(P0V��%*�1=';�y�p��%�d�U5�	�C?�W�3��6��7�.��؜�F��l�QR�T�Jag;Zӆ������|_SkǅS���JBV%�K����"WL{���������3%��|��.�v��,֤���Rg��S��	�yVc��P��Ƨ�WRe%O���Ԫ�7B��Q������5Y�����2ʞ�^a]�n_)%a����ɤv��I��5����m��j�YwS�@���n#�l���Â���`�6Jq�~cѨ��ȝo����,J��a`��'[[ķs����)���Fl�j2C�mתו���L���J<g&���g(�X���Ϯ��^�]۝�5��^`���$7���,f呔w�F��0KvE���X����ͦ� �ke4��n��'�{����ۄ���ӎ�-dᖸ5c�:��|�,���w���k����U��m?��V��K��(��zx��?A{vt�3�%}Ѥ�3W\�l�����M9���ٝFX䨗����2>�L}	���u�c���c���T�FO�����[+�&\ � ��>@{�"���y$�	���)Ž�����G9�1x�=.޵�9���	<�vo�U}��9/S�����i�!�yHYM糾Ox5�A
A��E����x#�oM�Eb���uL�wj���笠4^?�Q���eT|�A�G���:�ޫҒH.��~4̏k?%m���u�U:�u`���H뫣3��ͯ�Z�Oo?�>_T�y?#taT�e�D��od79@�AU�v���\}�EK%�n&ڎ��K�2��;vm��g���A�n�#���A4^\Dhx�R��Ւ���g��Km��Q�΄�^��y�x���V����$j�\��.�ћ��G��2_4UVd�54w+>��W�Nv�_����<6��������7d�ٝ ����b5���\J��z��Po�9F.���V�P"s���x|㩟���Քg�ri��)�B�^O�g�_����#y��ۖoЕ)�h��}�J�)c�Db��b���t�hU/��OnfsC#�ZjZ��;��̦.��>/�U�D��8�F��U" j�3Y7m�1o^=J��ׯ�xs�L�D���"�!3|˷z�NjѺ?C�p���ZZ;�~�[��"r<���*|+#Nx˄�L�O��u����LPѢ���v|��?{2Df���2- m�G�\DQ��ok`ա�ʯ�Dc�Z|ь�^#�m>u|���Gb��q�_��|$ꩅ>XK{�I��㵣�$�/6�$ۖ��0�K=I��q3Z�g��2A��J����Sg�|�w��IT�A䈐� ��w�]����c��űO�?`�z`64��sVE)>Cʭb���a�ԟG�>�|�h���5�N�vLu�o��i�~yR��bDN^l^vmD��F}@�+�Z�x���I�@ԙ��� ���a�zb��Py|����Z�x@���[�wO����H8�e�^b]��b(��5"�R��]ux|{v�&?J�������^G���_Ӏ�F�q����vP�r|ٴ哀l	D��6��
0��b9��3ͱo�b��P��04^�h����P�����_i�"
��aH�:���~�)�4� �d�C�t8R��<�f�#�q@J�0�{�����
,��Uj�����Xph~
�^2��S��2�o)�ѩ�{2�!��D������>eYXğ�>�D�>,h�̂~A��V#dq�Mh�hK@B�w���v摒|:_��5CE��>�m;�M#�3K�U��AܞR@����B?�����+�(��
��笊��4V��G����DɄO�����OʯVˁ�LH������kZ�עmِ{q|V�<�R�%�%Ҷ@[�+�����M�H�(;���wGZN?�D�l��
�z��$�7czEyw:wl+�/�������m��#�_�g�a��9��]���@ꨌ?̭�"	q��
:j�h-C�DE��� u|�Z(,7|X����T��&�����������y�i6��ޖ�]��|WY�,�^�N�
�s)��`��xT�(�"��k��L��R`m�;M}٩����G%c+K���Tz����,��X������ǎ�i���]gMTYt�5��Q6�J�/�Z�t{ʰ��7��e�j����E�P��y�S-�ܧ�Ʀ�����Bi����
�׍6���V�m� �:�[H�d�1��6�D}ѐ��gA�O�ړ�Z�JF�?@��	�E&��4y�9R0�(��&�M#^fgX�5��!s
\�?�L�����ߍ1g)H���3�L��F����R�m�_LM��#\ O)�ڄ����mWVp+`�ߐvn�*UO��L��gD�X$!�õ�G�j��c�i��9]4O7i8�/��5M�]� &�Y����*��z�'��W�l^���I{�0�E�t���2%Ҷ{�b�f��G���r�
��\e�B�%~���Z�ax�Rg���&u`�|���%���~��x4H;�g���vB�C�UT�ج,�._#z>�*�m�/0=���QY��&#n�F5���`��}$t�s���7��F��e�b�TקB8(��Fg��@�(�)8�4-��
%;����ˌ�?7]H��@+���,���Cpwv�����m�В7.*�y��q�6��ؔ�藉�J�p��M�V�)x�n`�F�IZ'�]�?/�	�V1ԝC�� ݧ�F|�B���F����[A�l47�˽&���w�Sc�[��Smx���<��\�uJ��9���t�y�2����#�[wP)A����N��)���"���&.��#��iz���`�dv��%�'�ئ$��jC�cQ�f����l�m��(0�n�/7GS�K�d޵���0�F8EbP�����-�	��+?I�p7�@�fO����d�5K��ð`��v�D�cK��<fVN,a��=#Q�����seN*����R5���@��L�N���'	l̋��g�V�JU��i�/[A�_��H�K�-�3ּ�Vq�!�h���C޷&�y�W��*	]������72'YG�+y6Y���*��"�W6~��7k�b�z�M7�(�a|�uv]z#����Ǚ`��f&�����`Xⴧh���R��.���ň
�s�:�.� �:��%��m5����۔�qk�ʒ(�%n��;ҷ�\�F:]�������jϠ�=*��[��A,�J��8�Ð��[���Hc_S9h'<�_�)Eӂc�02�ŏdR{�vW�a7=���� �~��!�e=T�	5��7����3�¿�����#&�|��W~�G
�ZӢ�h3��@�C�vJ]]���E�{�����y�LFM>	��y�N0��m�/�Ħ������rX�c�~	s~5�{L|u�P|P�C���z��o�D���Z�����<��2+ZK�h�0Ȟ�*��� ����g"ъ��bh�����AbYX�R�qJ�,mt�`9�f;��y���N��%!X��.cXq� ��\��'q!Ѐ�x6H*y9���#��%l�^o?�E��3�:l.�l�[�ȿ��V�*�h|y�����������[>���!���^�Nsz<����X���WK�nB�,%(}b�%~�K�!�95��.�{� ���}��prG^�e`t�6�˯�{,�r��?��q��^��,�8�t�ޑ���e�_���9�)�n�*�K�%�����+��ᐮt�ֵ�_Y����L}���8)Ǚ��FZ""���6=�m�
RK�ݍ#�̷��B`gAknZ��Ú$$5�m��Lhn�}X��`�e5����O-8�NOV�����×d�嬪��R��M��K���^�D����;Q�+̐����{��U���?�Ǒ�F6����8~'��N����q��^io�|��XG��kۆ!P�uP���n}���辺F���{��/=Y�j��(��r!3��o��ד�����<�K�9b\6�-����t�y��@FPlg�Cm%�#��OI���w$����qPh�JN:'���W����`Pi��܍3�Dj�g���{[��R�W��>�eqFɗ$R��\�5���,�z��>^�}�xSj)���ۃ�U')=6�"���RNa����#�B���4�Ugf	���H[)V^����-��n���r`�ltٲ�m��Y0nOr2C�n9���n��em-0.��V��kѼ��[Z�.� ��c��1�a�Vb��7ڗ�������KI�ks�iN�M�D�PR-���Е��Ȓ�F'PQ����"���S`��x��ZA������e繦t��d3��_�i� DHe,�Nss.�����b\�$�5�Ϯ���M�x,����29�T����y��ړ�ש����j��	�x���vg5?��{�nk�lb�EKߑ�̩�+�����,3��ZZ}��%d�פ���0&��L3��|,��ɳ��_	�}C���Shx ��'�솃����j��E(]jM6+{ٔ\uP����[,�֟��? v�-�ל�`��d�M��HUƤ�p6l :0�ْG��#�!ZhiV[�C�O�+�>�{}���zK��n7����>6�?M�U.r�Uj�/䌴�����U�b���J�F��v�C���!%8�<o$�:�E�3�9�vD�d�!X^4�_��΁J|�w&.U��Im�iz!?�\:E�&4�L,R��ǱG�0P��6sQi`���oӉ]���hHn�:S\f���a��K�v��n�d�5q�_lC>�(Xx��@T%(�����`�e&�CR˺l�6��g|�LnU��+��3v�J� �1B�o��Yn�6o+��^��0����ൊ�^ ���0��s	X�rC��;h��N��ԛ��X�Ds�8��#�pb���.���9��]I�Ȓ�u:0S�)|��O�	,/����1�E�,f����1���_m����$��t�=!��V� (�j�}KEb�I�@�P�^f4�IhӔ���gd�������|6�� ���&uH:a�~H3)B��b�v�ͨc�z��&B:��b�NkS�e�_�J�C��\�����V��"�=�a}2�q������T`��<d14�e6C=�C&�E=dG�j����}���4���Y޴�)���KjD`���Ĩ�*�;�tc4�(���;\T���НLE��'�
n��s����s#�d3 �������8�S�9|�F��'��%'@TA��x=�����10�'���6!8XF��j46�ݖ@��)մ���S��h��n86��Y �U��R�����a�����T��!���M���㇞�1�+:�P��쭱v�͋xؿP����(�����Y�0c��2�R�=W��i2�7��͗��L��:�P� |<W�w��l�9�Ζ��-��}u�93J�ߨ���>ni�����E�k�nY*8M������\D�S*�ҏ�wtdNl�r��e�BU�^�^�.�_���	|��{��o���R+�L�n}��:�5��;'_JuF��?>�Dz!�C�_���݉ף�5Kե�Uz������"�w��z��٘g��9�c�Е�h��7|'I��vs�e�����E-��/������E�J{�C���=�I|qua��i-�^1��pk��Ȏ�[TM����8��6f�~ʤ½bk��R]����ap-<�����vr9sh�*��Nm�:>�-	]#�!ȶ�)����*e�ǂ�n����F����E��ԡݸ�,ˢ��>댑��lQ��lo/���ԃ����	Ϋ���;F�'��m�.�
��f�?9��n��ꕴ*v��Gh����ޅ	dG�	��7�����K<���5����\d�e�g�փ/ّi��R<�Q2�-3P��6��8J�v�ֱz�N�A�k|�'E1Ւ�d�`׭��C4̆�ۭ��1�@�bI��;�n���C�4�s΢�s4�9��M۝Գf`N��t����i�_�o�:.�����f�2xܾ��E@kjehj��������dkO��>oFM��o��6��a~x�0��!0�[�6��{�K�����g��bF�=�n�	�l�nT���S+G"/�za����g����h�ů�>���B��O�=���(�B���G<;�(���"�y���N|Г���Hg�����w1{DS$���t-�8�Q+={ن�)Կ�tW*�)����ݡ�E¸=����}��p���
m�p�´�p&��?8j�+o��/`�ԛ��U0�|ZY�M7D9U0&=���a������k���Z΁6π�W\;*�ԉI2<��O����{�q��K"e�	G���AJ����(�@<Nf�&���'���+���]]�� ��Aٲ����KTp��<;8t��4&NZy�r���b���vY��ƺ��!b�Kv!途z��m��X��6�XP3t�=��`��v����q�j��¼�%��Pn>e��N�G8]�.��w�@U��ҍ�/e$��m�U�ފ�6j+P�n�65��74�%����}_�Dh[�ͧ���&�����E%��J-��j!^�rS�9ԙ�G+�k��5�KZ_3�6�횴�8�χ�,MV覒b$Q�4�9�Z�Vk:��=����%E�Ɓ%g�Mϖ�;��A{�4�����VY�ں�on�l�/��p|z����7��ٯ�6BV_v�c�	�Mc��W�"y}ţq��{�9�[�`�k��%R\!�Bw�A���W(����j��z*|]09Ф`��f>��ՁF	���n����y�=���t�W1�њqB��b'JHJP<3{�H@��^�)X1,��WU�߄>�u&1L�?���;R��ɨ8� ���qH�C����j ���=�M�=�(�5���*ͥ `nS|3��9�5B��0�`z�<���ON�f���@�y.���E�X	�U$�����&{=U������A#M������P��Iͩ:��Wa�6n�(������ht����4:�G3��UX�F"Z w��}4�~y#v3�k�����2��L������#����ԁV�+:���]d���k�L3^츚6i�j+�۴9J������n�I�>�%�.(6�1,M$���"1_j0�AiO�J���ґ�`�[���d#VLC�ݶ�cZ%������w�ƭ�fA�eW�As������[�2B���c�]��Z�6Z�Ғ�hJ�p[$S �p�BF𩸉.t��O1���*����=���4"y;�C�!)IfE�[_U6�)f�����[��F]v�����-U8�mp�ƼS�������~`�l����*-鳹.r��s��,`��$g{��Cj�NU8�>H����7� m�`!�i�*2'o#M�C=Ιg����Ǆ�3�ϗ��:n1=�|����a �~�v�����,X!/\ҥ��� ��[q�娽.�0EW�;G[-i�+8�-�kxQ}sJy@/	$!��ZYџS��nY}�!�U��d�w�Rlఋc���n���G$Z���{uoƹ������2S�J�E�g������D�MU��#��B�""����I ��c]�H�Rw�>��K6�Hd��
IRHi�b���i��藈ic_�Z������!�|3m��@G�1�D��05K;|�SO1��Ͽ?JF0"�����Wӱ}��'�a6ݐ`�T'��AiRnX)����B�L�B\�J�6���8�Rc�x�ˣ���+J��1'�̶t�(9�����<�}W:�t�,�Gbv��Ri�	V�x̵���`��E$����=Cd|	dS����B�w.�i�3����Ki"Eψ
5�¤R��<&����5��N1�����f���K�m[z����ry	�Y�ZsIdS��PxM��i^��|��]h1v��K��,v�א|t]	�3��|2��\2��DG1W�������_[��z��BB|j��3��]�� D1L�|Ɇf�q�W�h��a��E��2���D��ӈ$�6,��>C� ���a�|<�Bt�����4	&���Z'��.�zG;���V�pǶ��>��`M�������� ��1�9�����Ӈ��A�`��Y.+��х�t�2sb��Kn-(�w�|-N�����s-0�*R!�'f�"<�G#��D�-�]�&��	�!�$�a����k�j H�Cݵ��qY}�ƈp�w{����xI��ψ�>�یt��+8WTZ���^����H��]�����$����Za��GWWPȤ�2�����%=27{Qy�%�"�`�T�s�N�ϭ��٢k3�����I\KvG>��eպ�d�Q�^��D/�$��^�o�궋��*�^��wա���>[NC���e�����=�l.�K]5��T66�ݦ��e��ҽ~=D��&�M��Sb�����oę��y(�G>�*��<u��ӣƅ�E�Sˍ L�4�����Kh�o�������I$B1��וj\�>��Ǎ�!y�~X�6�m��~�xA^vZ��?`)�7�UY�H�-�:J�hg	뗄�"L�h�<8M-��P��;oٮ3)3�J���[��݀x,&����h���"tک��N���'�7a�;�p>�I6�x��Ƀ�VJ[5L�M���٢V.���}�\�cX����
$���}
@�=��am�/	���©Ce��%�J���F;�ǳČ�v���ܛJtř���Ȭ-!<y�|_-D�~���xA�4��h�n�:o�"�A+U�2_��>������忁�t������X��(gq�@�=n!���D�^�N��fIK����D�2�'sw�Y�t�U��5L�?x2�z�ɝ� 3\���[�����i#���=���0h���q��ߥ����O`B4H�8��_Y�������\݅NV��M��ػ:�A��R�`!92��ݠ���Mp�i�k���m��x-X^^~�g�;�'�;5��"i��9c�.�3���/��A?2�֙�ԒڄDS@����mQ�m�/�9t�J^Se��-|�?��_Ǉ*�{���0�v� Qtl8�.�ܡӼ�jF�5��5{�ܝ&f[֝�ҙm��K� ��~�h>�k9�	�XImo�s��w�^��5H���t���k^����D�6�wJ��� ���0F�mqX����!�\�8?;|D�����kL�y�d3�UYs[�YVy��v��5��W�F�4A;b����\W�ak���^H�pj :�12p�b�١�S�����d�jG�Ys��ϷG(��ڍL:�oo]��Y��c;�w�WP%�)�?K{�T}��������學0z=I�6��o�P��l+.��ɀdh�{���2�����=%A�"��%�
0������j&����r�ҩ�(���?�����n�J0�q��V-���-6Nӆ��^9��`�o���m�ZKM����I�a߭4�ϲ�+�f0d$�	W��SP�c�5:�c�0f$���,�k��Z�V\�y��읆p����W�����z��0cSB�k����xBB �����'����(�GMA~b ��g_�&[��8�������H���^TD��y�tS�Q�s,\�1�6�nQ�kg?f�qOѱ���-��F��
iR�Yg�"��%d��m��@t\�v�lnh {�y)+���E,���Z��;�~�w��M(գ�i��鲚��E�*鍂$�Π6��9����s����v屷r��1x�R�(�R���nZH
�^Z!x� �Z����W�('�/��r)[��n�ۄ,)����^y�j76��x�^}}_�_B�E��>}@�ب�f|,�	���_�ϰ�ۅG�#�6$�(�Ev�������Y�E�~�j�s�l��][Nv�n��G�/߫E\]�)y��~Q��d^智m�S[�U�o���������pW�WȺv��-v3� �XW��rzKdE�'��c-�HtH5�Hw.�/r� ���T�!n@7��ް�hs2)@��K��(��Pf����O��+4�;Qo
�(�G-�������nӚ��m�U~�>0*-¿������D�ym��ph[����M��󦹵 ��Lv�;8��p���۽������!o���f���ҫ���c\Z�A����h��
��_R*\;w�����;�/N�B�x��ri�4(O��^�W�g�-z�3�fH�X$�Eٌ��yg79s��ӱm�UM�Oc�6�Ɨw�,�]1bh`WR+�Ƙ��c�]��ο������d9��Qh�34��Ȟ�>���bC�=B�+�-�f(n�D��V���+m(3>� s�:��=�������:x }Ñ�I�}�W��/�/���_�����6V�ur�twJl��+�!bN`��M�c9m�dI[���}��_mQ���%Lǋ���~�_�4�:=�������Oo��p��V�+T`��S4��n4Þ��x��^9>Ǽ|4�*(�#\Gw���q^�"��9���M�8��6�����؉Ij !��ʌ���D�a]���!	�ر�J`0�ʖ�fˮn~C�P�j����Z���y��qA[��1}s�C�/?ǁ@��Ĩ|I�y҅_\7?a�CX��#S��m(��'
��y��~�?��8�h׋��0=H�f��@����1����Ex�J�>p��'v�n6���T�+��)wA톗�����������h��99�B�ԬW~/�:�e�G��i6Ue�<��U�6���'ڂ�j!��! "�W�D.�� b<��RY ���Elŗϛ�֟�T7,��LB��eN���r(��x_���Z�~-��%��Zw#�K�,�Zl$�i@ip|�e2��_��	��+���J뫉�*��K�Z���}:�E%Ǡ���=�9o��A���zۼ8F��o��%���N2�)�7˒�F��*�����|KAj�uV��`��n��!�O'|ٿ�^��V�n��+]f�n�n�~X����N^]� �}i$Pԫ
����B�6��PŴBzd���`�:�[H�/?� �poLP��B���E�m��|�ϼRT9E~�_�	��o<a�B��D�ԛ3��v)����ڵ��9nN�&�4�o�:��s���.�
H'KQ�-�y�?CNX�n�=Q�c.ȚK�8˴�y���*8b������j�ҷou3p���vN��
��6߾h�:�5��h�D�1�d6�C���$l׺)1ŸF��%�h0.>�
{��L6	���\��hr��B����13�ߢ�AI<�ұ����ϰ��2K������&��y��g|����ǥ�`�BFP?�C�u��AL"S7lp��B��m���mcJa{��ry?�)>��A�7Bf�M�����ODӮ��w�ڨ���B���7`ݘ4:I�l8#̐���5k���y�샅������"��$�PO�$� ����~Y��f!���cp�4ԋ{�*�������F�J�0dp#�pF�1/:�:�J-�z��%n�|�ի�-HXTa�K��g�_�]�x��e4�S0���5�����ˠW��:�����)1���_�]O��2	0Z�c!�;�Qq��)���9�l8Rk��|�-��>{�9깎4�^T�v֙�\�	����wmu>�y��c"��m������t�/h�{}]�Qx���)��G����H�@zU�n�u^����u(���[]Z����ɎǙ$d�Т��k�<��W)�����ܹ٣&2J���j������>�����7�:T�Js�C��C���5S�7��x@�U���R���7���^A�N��|������+'H[��S>$�'����s֋�d���-�1+�_P��~vk��&���soz���2Ρ����!sm�A���[�����w�����w��A���t�af-�E�O�l�}��Z�F�����M[��8m��J�"�܁��:�r؉j�'^��t-��R���`��'L�lk�:]��:�����4 ɩ$E�/��dZa�3/����'>�$��C�d_D�I���)>j���d�A���X�)rV�J�a�6���:I�����8��+�-X�r�9�I�qz�������a6�tDh�J#ab*2���2/�ٺ��5�nH��)%0��d�ĩ#�7`��AsT�q�b�G��u��3�3��ĤΔ��)aG$;9�5)����_�/�V�d�K�;����u�؏yPh*�:��:xl��ok�y�l^`UT-�Hԫ$��Sy}�n�)����I�K�Rn��+G8'�Z锆�	�	���[fS�墾c$XBz�l�,�`���O)�Kd8u.G� �0I��U���@�Xx����01�b=�̆��2E�ѳ�{?}��΁�7ϧ��;Շr �WԡU8Iyo�5�

��(&�ș�U��Z�:=����2�u��O�;�v�&�.';I�6��]m�]�M��]!X�ؕ�"G�]̳ߤe�w-m"�蓗�c��ؿ�Jvo�[ﱏ�Ǩ�mB�F���!
������}o��J�,*�*g)�ʹ�_�f>�B���N����(����ؾ��_2����V��ha���i[��$��or{�x� �Ⱡ���a��hA-��m����R-
�����<N�˘�\�`K����Q<��Y�H2 �9�0OL�gPxh����K��KO��J�9��7���[��9�SP*��=#��Q>�������Iy��wo�,pw��aܼ��=��a`*zZ;�����N\��9GN�>��8f��;�^C2ߞ��_L'��G]7w�{��r/M�[���R�$�.i� UP�lX������7t�1�Ѭ�v�u�]#aRl�]1��:L0�ա��V7���#(wp6�bH�J���][!kI ���%�ED�H��݈�y��f֥칆V���w��ľe�r�Y#wa'	d��en-�s���)oq��K�J�Xa�#��L�����81���+�Yʣ�k�$���N1�� XS�s\�~�a���YfkKPa/��.���1�����H�[���م�����x��;��P�hpg��#'(�5���?ڽLp���X�_"�&����0s�D�������H�k�"U��`���΢ѩ��c�8��_�a��x�Ҏ�8��¾��������.5��(�eac�q"��X�`猿O���*o(�#��i&���Z�܉��/������ \�:��<7Ԕ��.Tz[�0�R� �YG�b�G�V�DT��'��Z2�(̕� ���{���5�`<��͑�H�A�7t�n���D�I������
��s'{���H�S$�?w�X+g+1�	�,����V�b�x�@�vg���ˊtC�W��������?	L��8��4_7��8��)M���AS���M@���<.�e-��^3�V�����;���#�}�X^�Y�����Rb�{w�6O����g�{ޮsb8Z	�xg�/(�)Y��!9Gk�����#~��`yj{�?�bg�)ha!WR��e��2��9��H�Y�.B�h�!�����͔(������`�����6�> _�%��v�k���&�����DP��߬�q�w����";�����)	�����~])����u�↿a���j���AO��Mڿ�H|=�5zoUe���oD��q� if��k,�*�3�H�N�������LJX&�������-0�^M�l����JK�^]�x����2�C��H(�]����ᵛ΢N!6�?0�u�;@o����O�XBo=�e�K����[C`�,���N ��z����da�>��QP�>���J��A����HBk����?�03/ЏD����8�W��ED�#���ĤK{��-�|,���?������J�-��%���?�o��uGӧ��Ȩ�ǯ��1�����ˆ}8B�,���ӕм�c�it�J{E����7Y/��nր\�?�SlHf�H��q��LOdy0����'�mP�a1~	&J�y�?����̜�}��be,��j=-ݼ��"��I�#�����0�. ��Uʐ�K��Mz��:9Zb�N��8'Y�܁/R��G��+?a�D�����K���{�*e�`�<!�&M����iL=U=�*��ՂGr�q[�]�G(D��f;���4t����*e�*��;q揁D%	��C��uYv���V�l���Kd�����z6��k�h<�α���qE)�Z_��q徙h+$ڊ�u��
��]<�� ;!��"1� �����6��P��ɞ�/H}8�w�2��F�y���fvܧ[�9f.��(NT�|�j��~F!�B;�s���r�'�g�O(�֓��jz�����k�to5�=9t��i��vN\6I{{��6��i+���Oe�����9�ӽ�h��J�#�n��U=���&��:ty��n��.�<�{�}�b�r �MC��&�����6ZCa��{����:b�����0�T/��1�l�¦����)g�]Xē_"�J~!)��v�I���No��˯n���ΰ'������OEM�� j�ї�s(��v�����j��J��*�u|R��1ڟB']����}:���%�}���3J�u:y^�0�J}��$I�����`�!U�P�d�"�t�*�h�A�2X
	��C�\��ڡ�\�=�����Z�ҡ�q�mn9�����urňr&Yp��H�wGO���&6{�k�˔����.���5�L	��Ij�6���Gm��c�*J�o;���֛?:��}��c��ݞgs㶷�݇}!����N���3����#����������X$ϣ�����K��]�湺�ߞLѿ����|ƹ���%�b�������%I;(��
��\�u����X-��e]��%Ǹ��F�⛉o6�|�}l c^m���h�rT9�V�K���a�m���4Ց�,�oeEW�3o�gc���J27߹PW|ډ��ߣ]�;lNp�v��Hie�Fy?l-�Q��� ����	����mvչr3>�a�����2��`5�3�,U��1w}W�]+�RT�_5W'��W�����$�� ��Zh��l�v����S�|me�D:|S�)�kX܀l�h���VKƦ\�7���w�l�:6�X��Ab?�ʤ8����-��^BD�.Dv���O��J9v�"�"!4�#�jU�Dtv�V[������l
܎�J�u��|q���HW�ƅר�y��֜���q��t�9k�`�F�o�5 �$n��ر:SA�m|����\����A��ݙ�i��]$�8��(��27�R�2Zz_f���Q��f#���?T�J�,�m�f�~�f���#���%�e��J���������ČzmVxe�o�"{�R�K�^�p��fg���KGo5�33Kj֩��T'Q=�һ4Xj6Z�X�a���]�;���m�T��SD4���������o�3t���|��gQ-�`ib��Oɓ��i�w�!�=tT��ފ�K	 a�ۘ	\��Y&���SL��k�b��h��J5Th�7[�a>9H��*�t#��|�_4d_g5���%QM������φ�!UI
2W���D�(���Ю�{�3�t������3�%%^T����������t���'�jܪ^�y�W%h��>s@}[@"�{8h�'���V]d�S��mͥ����Z�#H��^��nG(u�� �}�9�`d��#ܾZ|7����\�!CG!����}��>F[
�Z�T�$�M�`�3����Coo�i������ѤT�~��y���P�k[�#/��� �Uz��]ҧ6��&j=�ߚ���Z��_7�B�Lc���U�7xo���ۨ�k��ӎ]V�i��w�n`�h
�kE��O�澬�k|+�I��YG"�|"'�F��,$��3Gh�:��-��Nr��cZv��q����M��C�Ʃ�˘�ʼ��=�]A�ǰ;�g��q�+RdF�sx�5�꒩��,+�eo�S�<O�+��<+����5�T�<z>�&Y��*q|Ғu���s��imq7��ZoQ0 h�GW@�JG� "r܏�V�è�ٵ#�\9�f
"j����s���a ��+�@�!K7Z�S8�����W2��yȄ�HP��-t����]��ܻxdgstnp�?w�u ��FM+2c���E2�]T�U�����wI/i��&L��yKip�!�&Q�{s,���9�'P�*�����������JaT��=t��?���0��}2r4��S7�}�T����k^�{\��Cry��堩l�H�З�F?��d���Ɩ� ��`Y�5��սgr>�1���^�����Zp�)�1�g��W��'����W���%��{�njl��-����0��v�Ê$�|m#U��UE�ػb継#��'��_Q0��4|eT\M�-� ��L���������w����0���ww�3��Z�יuz��K����9��8�y�O���v���כ��K�s��]����تh7$rP��N;�L�׃O��S���
��Ϫ\�96�}2�\v��MR��P\���ݷ�=�=�]���Jz��(
>y���.Q���.�'c�Wg�i�h�S�� �t=����-^�P:+{}����HYB�.�6�������DT-��o�|M<��`��o��̷VԻ�������OO'V��6��HU���&h��>׽'b��)AJ��938nY�<�b<��N���8�[+������Gx��놮��FWL���<�)&V>k(���mh��_/ f�����;����}2�C/;���au(5BAVs��m���ꍈ��~�I󞰹lb�5۳���'<w�g����m�If̉����3,������'�<k
h�uZ���0�����V��������]o债�;mC�-�`��� ���&PY�J���,�Ͻ8@��'����4�7����w�sl� ���g��:`�-����:�]i����7k�k. ^���G`�W��y]@`%���uLX� P ��	�4Ce��û�!类�H�f7Av� v1z*��WN���v�`+��y�* ��6�^f�,"�#h.��ǰ?WP����&�v�^����2�����͓c<���d�_I��������Q��bEKkv�*�/�<n�(s�l�e����wT�h�^T��������$�}���I2����zf�ksg:6dL�-X��;<ld�{��s����e���j��	��q���n��O�%����8��ܡ�䝈� S9z�8���ô��2� }���
*V˵"o�ыr�2��_º**�]2k���8�D�v]<�����F����+���{�U�V(�	�6����8A�A�r�]��n37�PG"�h�!�8��ݸ��y��� ["�?w��@Zթ�ʟ*�5���� ^z����g���C�t������)��G�$�e����Y�ev-]yK��H�͉�����&XkW��WՎ��`Dg$��^OW�H)3տq��=�.�K�qO��09	M��c\N��`0��TL$�K�T���\������&��r?���x9YM���44�biG�:ۦz���x�D��!~0�Q��Vo�7����`��l�+oӭ�R;���AH̳2=F��ШD;�hx���#��ۼnlM(r��ނ�
3���a�����Zn�����^���O��|��}L�h�Z5:�JJ? �-��d� �B�����ê���N���}���n��m{j(�8)}cGYP-�J:e2H?6v�T�W�G�&n�m��ya�V�@��Ǆ�$�S\0�ܹ
��<X�8?|�"�
n����NOZ�<��u��F�9�?#E�����O���"�K��`�)�%��e���@�#��~��I2eԤ:1�T����к��j��c5��֧�x��N�8)g�(^0 @�I.o��jғѴR�fx���u��QSu�~�5e�n�������e�*C������k+��P)/�9��K0�����P

�e�&x<q�7���a���O����G��Җ��#._ٿ�07v����� �ώ���gA����YU�ߧZ�K.��D�Xg6S�L��k��s8��|�N�D��C�~Q<o��9��^|C�G-��UʆW��m��J�Qsɱ�¥�~�m������+{8�����0s��[^g�I2W�e��<kFv�L�ڒ��5�n�^�*�.�P]���������/��<�_�{�C��;��U{n�h�?˒�dn��R	s< ����8:^�C��Y�h�7�=$���Ӂ���	�ڰ$���:�-}�jJ�c2��^Z��)�V�4�C�\g9��79�]�=��q�|��������։0��S��䩮	��J|,t����8�J:��A���aD+vvZӝ��kH���_;��ӟ%�M9
D5��嗑jQnk�퓄5�2��I�.	�Eok�,]�C�Z�v��l�����( ��<���kBA�/��91<]����[ѩʌ��+(C���N'�&��%�%x����Jxn����3jp8>�4Oے+L����ߏA6�:U�%�SKwT�ב�M�>w�,@����b[
�&<�s�!W�����Q���M����j��g�g'r�@Y$��ď���[@��8�<W��W��ȝ�1i>�V��>�Z��\{�98�,νƹ[n�yd��HS�����4����GK��R�mR���]�=�<9��a���.'|kD*�>��)D2��f=����B$#�х���Ӗؐ�L���ׯ�Pԙ/�ȩ10��6W��Z��vC�0<�UX��x6z�C��h�JYf�\��/O��z�F���F���yĈY��"��'H���H������N���C3}��@��ibn�.����*]�MX	P���~�ʉ�kj�R��z��E��A �Y:>>r�ɉh~���w�{�a����?*hO��/��8�w�`>�����z
#�ԝ�R]2je\/Si�KA0h[3��T�� �W��k�|���FG��a�����zS M�1���zJQ�+��̹"�z�%��M��0>3�\a�MY�����<���o^Ǒ^�gV/B�.h�s�=��<U��f|� y�0)�0�&��L���G32���RR«��Us������D�FL<���M�б�h�w0A-ҵ�[u�
gp�ļE��A�K�,dn2�C����Ne�j�5jG/H�T��Ԓ�r~��^� �|&�&���T��L����X-�\*��Z$q�iEMq�]q~R�N2�b���Fv$ _&�C�C�Tcy~�6�Ή�� T��� �X-�l��n�^��d��b������&�bg���GF��ݹ;t��	޾�xn��������`�_1���?"�\ؤv��dk��F��Ѧ�t���)�ł��yu�?�`̢����7k��Z�ň2"�~ʭ��j�h��z�_�]B,%�[���+6I��LK{��^vi�Z�)cvX�FP3��ֱ�=ଜ(k�l�g�:�L�h�i�ވ�	ʯ1���e�����]��4v����ᩩ%>.�!��܊
�z�����xL�o-C�.w�����~�����yR�T�݈ݏ����j�2[y��"��XU�Iܰh���ǰ��3͎�E���	��nL�g�4�+���y�6f����;���"好��)�|�~٩]0�ϸ��d�F�)6;�Y��*v�ഹ檧�c�y����}�cj{�}���(�g3�O�������+(+._�&��kfzگ��(��f�)�@-R���KLc�8��ߓ�w�6�}�LaR� �-+CEi���D���ͺj����W�Ga�5A�n`'g����"Ŋ�����V�W�Jr.R�B`H�|`*����涔ک�) �$g2��c*�?�H�kYY3��h,$�FP'N^K+2��4����z�Z�� ���Mo���f-�6\W� ��"��َ�X�Q�s]
p�3�� ۸ ���os;�np����Z��4��Y��'M��9�&Jjmz{�ʺ"R��>�'Y߬^*�����pK_.��+�fk�#S+�tlZ�̧SsվSb�2�{�ea������^��\���c}�c�@���Ӽ0,�S|, Oy~~��f��ֶ��}{{��w2薻�nNJqt�.�B�q����X+�E��%���9��y�6^)���y�D�6����Ԏ?^���k��	pƩ�s�����?��[��Nb�wRk�1��)��4ݻ;������M+�x
����_�UOu��@Ax�4߿M)M	%v�ޫ�qo%~�ݐ��s5�}�1���T�%���f�< pG�[P�ioo/���ܻ[�Ɔ����I�g����f-�t�9k�7	�n�k�^)5��F�fc;��!��u��1�Ic�//=��Sl���>Z�u�
�O�Y0-�p�=��Ɇ�#KZ� I�$m_��{��Q�cK(�m�!jwk-8���0�C��K�М�#����_5��7�a�7z��7>���8�l
،Z�Ch��M]&o�Уʶ�0��e:=rI���@mgp�i!�pE ����~��]`e�.Ƒ�EEM��r�D���*-mj6ȃ��o����,�ʡ������e>�j�e���jl������ԝ��*U6��&�)��Ө�d'���kb��Y�"p� �N���/,=)TXn����h��
ܼ*�ɝ���_i�Ͼ�f_vs ^�B1oL�C#����������4sED�<�m��N;
�p�l��ʳ%D�s/]���L�DJrIccrK����nIj���)&	^�E<$k�&a��J2,���p��]w�G�����	�D?N��m<��'cͷJ޲�<5�c�^�
a=��W��S�2/�oT�<|n	��x"J�i�n���Т�&fXG��P�}��5J=�2����h�vZ�0`"�gf�.-�a��	���}wW�~��������Q͊�+)�8����՞v7n��np�^|ķ#q����M ��%H���W� h� �9��ED�����R���W=)��>v�of �Q�w��s�umN�t��
S�r4�*#H3���Ԕ6.���J	���z�
sx���^�b��ܞ�d�Ew���]�����]]|+�$ҙP�p�NB�,��&ˣX��Ʋ���x�� c����肬��M/[����bfn.���S�<X�/�H��΃�T'�v�y���2�ۅ��c����t��#���7��w4���lx����T�ũ�28��;~��Z�E*IXU��Xy?�`��yP�����S`#�%��FK�hy��Z("ӽ�kvv��
�v�������
iX%="�|����5����z��g��/�M�K �e�#�"��Kc �B�x��S�e�gl���o�@Al�L�6{DO��]CH~£[��@���oz)J���m-�a���xT���*����T$'��d�e��4<_�F�m\V�K� �`:_<�Y��8ܘT�� �����|�r�f���i��$d�$[N�O#��7n:
���Q#�`t�s�xJ�	|��&�eX)�T�?3�dS�pk��8T�?�i�7����#�L>� 
�'�M�����Tr㲭�#�T�i�,l��Cȥ����-��]��:J�zU5��=q��/Z8�'].���ץRE�~������aꗙ!Pkrr3h�G�뿎�Lɖ(T���#�{Dj�w9����I�`�e+?x�u2s>;��F-Z�{�:��AʆStn���UUM�5N��%ieԹ�T�.�(��mGس�t?��>a2��t�1��������ɧ���	�ث0*�-�O�E��Hb���Ɖ$��eC`�]�H0w�$�Fܹ�1���ʼt��sФ������@����̜�=إ���57wn�>4rc�����o��}����w�J�1�Y���Pm���mZ�U��y�QW�ԃ���TN0�������N�� X�a�� �䪤x�q���⫹�~��1�ېu�7n�I�^�%���jW�d����dG2���M��W��zx�9�~�ajJ���B12�n)l#���dË�N(
��_�'b�T+	� s�:C�ҁ9�{�`��J��TN�Q��m�jc��Ρ2�NWε���h�����(�f�}N����Wp��⦷�"�m�km
|XÆq�M�,{.
�ɉ����`u�-��Tn���N1,%%�˚߲��H�]Ȗ��n W���v�*���K|�RӪ�y���ü`&?��-�2����䜁��i� I����'ѶKq�p�1��7a�j����I]ɪ��{����������o�ԞW��������챊��e ���=��V�{Gg�r�\t���a)/c3��_Z��4ҩ	]�|QL�v�T#�:*��W�kL��D� ���v�C`��c��ܧZQ����C(�r[������Zn�:I�+�t3�"Fׇ��a����B�L��6�F�5j�1�ŝ��@�d���ؔ�c�Mg	���s�ϑ�v_��H˒�ڌ~�
�Yq$$ڿ��^XXȶ~,�&��j98�d�m��&�hqh7Y��􍊑Og�B�1�E��5��f[􎢼!�u|:m��Un3��h�B���E���\�}�@��AѾײ��訠/p�5ŧ]۫'0@	����$��@
D���<�nfs~>�D��\���N�3��<��"	rXd��2��_a*�ws3��Ύ��ŀF,���͆&��s§I� q�OP��7 F��ݘ�;����7(�]+Jc�_Ó��u{�$���j�b�x�s�[:_��?m�UV�T�I��v�*��Q��2���<��ԇ����J
�4(�~R!�<Q�{�T�O�����b>�����;(u�v�O��f<������Z+b�3-\�:N�O"BD�c:D�ْ�;���:�G����{�=�j����=�7)7���::D���v�������Z(��:�xo 茏iY�՗T��9ǉ���T��ja�����l�TLM��V�sN(��장�������G��Ѓ�J8��l�NC�#$�V�&�N�_��Bͩ��>�ñ'�c� 9`x+M�pH3��)�m���a>��ѩV��#��c��d�}M����&��D�N��N��[���)?S�~�%��N%���i('/f�X9��3�H�\I�݄��K�\��{�[w�Ȁ�LY~gZ��o�
����!P��H�`��[���^��{\�iA���V�IM�n���Wv{H䓷��3��`��3$���i�υQ/uZ�X"'�S�(}�@��F/�L��Q��՛���8? -E�ZDx�^��>nԄ���>I�o�~�t���4�u{®x�΀9m M��5���܈̓�[�J���nnk�>{!�Õ���M��'7����ux�NW�7UF�绐���{��**�����k�b�B���jV>~�;����A*��T[���3>��#�G�B,�v����l�+",�p������x�PiGA��8l��N�߰�jW-�՞2�V�r�mz���RQ~"�AR�<�^i؏��\�Q"�,O0���%at�)�hY�9��y��p����.9�D�Zh�ځ�0��g+����Ř�u,e�<�!b﫥m�2�7�o���q]��#���1��i��b�mu�w���3�m��Ә���?��1�� )t�D�g-O<�|��2��B�'�	m��k�O���@H*�#�mW{�NB��0����Tڻ��ר=�$�}|����r����Y� ��\�������΁�\��l��5�ȼp_�2(t�J;xK\��a���#}7`��Q�%S�X��.���.i�w�H*�\����A{�zaF��d���-��T������5-��~� T�s�n�]v����%�V|���,_7+����ݣ�g�����$V�%���J4B �"v	�᝺�i���� ��ĵ�j3���^KIh���߁�|���W�S�&h#nkL�:��[����,�`��>w�>�R<�5jx)J!b`a��v�PiR�2]��r����)c^}��SE(C���_/4׉�w��M���#��[_�������¼�1�랟j��f��)
���y��T�8��e�T>�]��4O�r)��Т_Q<���"��4L�����)^b�L{-I)Chӯx2St��>EqC����	v-�g�+u����'���ot�������	r�s���+Z<i�iL|�PF�0ӵ.�i��P�y������C�B��B ��"/�Ы�3���Q���o��쩌"��Mf�?��2������I*��
�;�1�6D�[iسĪ/��J$��6\���&�ی�n��x<�R��ʭ��l��˳zװ��IY�`�5QE�kY*=<��.�V��$o0�1�x3'���g�.O'1WT��b�c�ZQZ]����|��'%4����� �jv�c�B�'�ُ*��� f]U�.|C���H�]�E5��@�[;u��Q�c4D�Â��qpTo���L�*̙���o�M�ۭ��aߟK��2���z�d�V�Q���$�9l��?���
0����,y>�G8��Ovs����e�Z��9������yv�X1���bQC� ]g����Y+V����ʃg��/s'�?w�)a[�VT�h��x�$,�t�t���?�Bf��6��l�jp�����F�k�:��M+��l��g�Y�?�Hq1�9x���6������&Ҿkh�����dP�������孍�W�,_�I��6�p�<��p�|aa��~���S�]���o��y��7��-q�(�rZ��-�>�M��!�\�� ��RJ��V�VZ�����d��?��:�$r!����T<,��5Ȭ����12�K-!HǭK��-��lݎ_}�׋8����0ִ��.�b��c��H=s�l�J��-|��<��t;�D��#_B�s�Ҥ��QrW�� �ɐ�K��ܮg�a�ىɯPת;Ͽ+����Az{Y��j�&���9K63��NC��jߌ���V�1��u
�Z<��F�rU��0�)��z�i�"O�>[�cǥ��g�C}׉�Xa�tvŅb��WF����o9��S����r`{�~�)#M'�-��8�"����^�i�YfI��7�9Kσ�AUΝ�&�ǋ`�z���(o7 R��<'�LQF�bb���+�ꋪ�����jG���)��[?p��֪�j	잴Tַ�9E[�kŇ�?����N|c/�����>���Ĕ��0���L9d�w���x]���D�գ��ȳ��WxT��n�a��}�y����M*,m�moT"t�����pu�u��u=��Ծ���-�e��oI"��o+.c{��d�|v�
�0c+�%�v�Y�jIZ��}�i�M\ߴEܱ�;r1��K�]'� ��q�c.�u����y�X�;6�f���yLR>��ഋEKo�(��G����UJ?�H�E�ſ_�q ^�f�]zŋL�)p=�C��嫻�=���!"!b����m�>��1Ҋ��]i
�X��r�c��˓�yA�jS��'�U�Z
��Y*!V��=���� ٨���.~/�k6�̰G�D�}�zR�� �:CU%�@n����&�C�f�K��HA�_��p�e.E	��6S��!���̸۝��O|w
�@��T�,ǡ}��r�&L$�<����؅g
��:�{ťsR�;�ܦ��o|�w��Ԕ����
&GS'H�-�Wڇ��&o~�8I۫��1�O
�*6�KG�,���m5�����K��as��Ջ�;J3��)�r;���Ʃ&�]R|���4J�TE ��i�'�i�M
�M��$�@�"����NO��(�m�����42	o�X�L]�i���v�{�\$�O6��lb�^��#"�y�e<�}Qx���+�Z��^|u�4|�$�{��S'�����@	��	yq�u��B�a=,�X1P�St�f�#����qy�%�_�w_�7 $x8X�x]���r$���X��j���S���UU�Hi�jA�RJ�X�U+�H��po�^L��^2=��<���WN�e�t�
κ�O�n�1V��6��G��T>(J�t���3ݰ_m��)��eΛ��8&5T��A{�ޢy�A���?�\���9�2�>�T�Y�v�0^������@���5��ܭS��ٗ�F��X�j������Ƴ����W�ݟ*�|:#���?������'�A,Q�uL�b�J<	�|zSRM#$���8�}a��qhޭER\:'�L��B���`6I���f ��I��zZ�9O�^�<���N)[���ק �C%���o�8B��$	�q���|����Y��b �f67�V�P��"��7�<�	X�@�Z(ڄ��)��#�^�W���`'��O.l���1��Q���� ��������t0�&�Zk��b s��"3����[�����̎�u'��$4�_�Qt��Ư���,u�M�9b�ؾb�DxH�t��6��1���{���2�-��DB1k)��H���r�`\��*�@�ꜫǝ�-"y����I5
d�I4X-F=Z,^��x���:�R���Ƀ��ޥg�0_Ec�;@�u2sn��Hb;z��Pʾ4_dښb7D��8	E��E&M_^��p�����-lu���Y�;��H"ؠQ1T�J3LQ6D� �Tzx�lu���U�Ev�����٣��\ӿ-�M��X�	�Z�]P��x���{�G$�y SL���w�[�_*|����~��Ao;cS�>�X��p߼�/�_���C�Zߎ��cV�Oze����n���X&`}?��ڻ''��k9�$�0W(���C�/K�h$2�t�b賃��imS�P�b�������$H9��#h�o&���)��^{��+��&����ߝ^@z��1-v�8�[U:��*Jz�Y�����ThL��Q��)��c����f��k@5�pZ� 2��T���{=䢯�s��?Ɏ���i_���HBB�`h��0E��R(>�-�phI�6�&W�siԶ|-�l:I#mfUȈ�:@�.�;�MH&���s@�x�����C�҆���Μ\��a�Y�U�Um]�I��<���X���W%�1�FC%zM�"H����s�p�Α�y�j�7�����W�ݗ�E�r�1��/l���*L�Vc����w��K���s�x鯗��L��]_�"{=������[����w��E�o[(eͅ��Ć��9�.Sq���ÜB$�:��J��p�v}�[JT�P8#�b8��M��p. �p�y��]�|�y�w����B�n҆yg�+ݓ��'�"�IGߏ��&V9H\M򹛻Mw>𫩁a����k��B�i��M'� Ҕ� f��ix������KjL;�nN�;��J~;�>����m�]�-�aX� t֏f�©�85�_���-V����������Y��bi�/�TC��Z���N)k~|�e����79A��n�]1�4���:j`�!Uw�����tv�}�b�{a�ngi+�c0����P���Z���1Ŋ�iS�7o���/�v��l����vS��*^V��ΦYv@���6�:�16!�I	���j��O_VȕWܞ�WԜ��3��I*�1� YG�%�@��蒘���N�qɞ�)s� }i\H��bF�x=�1�6"�H/*Ͳ�?����xP���p�SI=��HSo<�7�-�p!m�r1K�<n�v�$bEw<�Y�\��g	L�v^��YsfA�q�BZ�D>�:�CƩ2v25�%�^��LD=�h�g��O�c����u�m�k	�*�t�����)'O�Kmk�q�T)vQ�{FQ� ]�M��&!fI5��zS �WxxD�[����r0�ZlQ3q���j�B�w�o8$u�\�&6Z�b_�&�!I�������9S�큣Q��`>h/s�.�j���0����.���E2h_VfaH����f1m��'[�W���������,��P s�"B�_�1�J2F}���x9���M��1��9�)����@LL��m�n�H�.K�LAѣԖ�6����mC����2j��UE	�����a��!U���<1���er�������h�)euZ�=r�M3��|��N�m���E`آ�A�k�nL�Q3�_g��Q5���'��Q�2N��
Ҷ-�1�����v�����]5�P/�xq��@���:��79�"#銡"MrSզ\-ϳF>���__L��h	B�7ۃ�2ѓT3�*}��RG�%Y�4YU��C����t��~@&fUs�
D2�6�:f.;���G���=ݓ�2��`�Qo������D�������;��a�ZƁ��F�_#4_��!E������_o*q����zr6�}g����"5��"	\�|-�P`[z��ڲ	v>�%*�+�T��^STM�NF�#�K.�=mӲ�T{��3&ҳۨϗ�������f�z]n~]�j��pd\� i$��%{�!�C��%˨�Y��U�<z����Y�0d����ʒ&�z0�eq�ǿ2覨�vW� ��Ic��H|<��W.�|�%�b	��^I,0�D��d��&�{��k3#}(!�:Ց��:��A�Ƃ���ͤ�'AO�t���B�/�ұ%��+���uqjO�¢��Q7vф`�Y��"a]�RP�Gn^��"��l�+�WsY2�#M��m���``�J.Og��w_y�̷��q��i��[��M��!n�1�x]��L�����c�k?���M��A���p�#�Sd�H��Mڏ�C+�jV ��D��i�P�U��X����]u�G-����j1�r=Z_��R��}���$`3�B2��g��KjNנ/�0FKn��;�m۫�yGNfx�m �����}b��0�i��D(ڙ ��;"���ץ�=כyaG�',E�I�)�`K���z%�7I�]<���'K��/kg�?�TК��f�I�1�M$K��6�w�h7�&�.a�#�)�tX�e�쫽I!���ǜ����>�-0��Xb��J��Ч��ԉ:+?Uט����ge�C���N��g����:$7rS���e���ʹR����o�V[������ l�S�r�&��=��d�/�nu������/O;-C����S�D�˗\h��[�����QNT���Ά����$sC�DsQ4J��O���~>�[�_�S��r�rby��z|�免D~�Z+M֧�?�%��G��^1xv��A�z-�\A���2�?��{XA��lp4��2��/�#�r$⢺$|����M��N�D�������N �D�>g��� L|���������h�!LҸ��JFw3��/��(fVJ9[�����L�t4y��9և���k���G��}�iζbUg��T8%��e$.i���<�s��-�oLX6@0�,!� ׉���$�!�U�	�t�����Ӭc=Y��<n�w�D�̟��W
r�pQ���!��?1���ew̌�z��!g�j(&�m;�O��bF��scc�*�F��k����gM���9 a�B`����m�]��`$)~�A���P����-�b���l.��UF�i/IK�x�I�2I���r�[&�l%���(1��P,���4�# �h��~ޫY�Z������~B����RĹ���%X����y�R��Y�}��a�M�7cn&�gةP=ě'���_ %���8'����WO�����sk�W�M#��(K&�s���O�X��L$��0�#_D����5��A��:�����]��c�����8��& g����zAh���1��r:C6�L���F5�jx����\����̷S��	�J�	����5����r�7�~�K>j��|����$�A�W�w��[m��COT{�E��Bg�%�V�;͔�>�a-���X�1k1�K��S���d�)��]����<J��`�FV`f�pv��p���e���T�ePH�+�w��K'��l_�뉃�Z�� i�} ���I�����4I�$d��>e�ڂyi������&<`0|�H�l?�	ΏBYP�[�JЖ�o�V�Z�O�u����A��?+�i^���}���$JƱc4]�U�b����K����%�[��)W�x���l�zf.ۙ�x���X�\~PP&������AY�r~�d��	���E��v(��P�ߢ� S9!�T#�4�ЮC=��<��C�Cw����-��8ķ��JCF��ɸb��,��`ұm�ڥ���|*�����nT��_�uj0�$+���ޒէ������&����EV�-��*ڌ:tV��m �� �$�i�^̅?'�^�Ǡ��cHt�{5�S,>�9���.	S�߰��?���%�t�U:W�o]�F������Rt�� Ab���.�ԯG6�'Tn%���������D[���|�Gc�n�pvU�$��Ĳ���2��������������8��b�������^)Σ�u��.��S��	g=���U+T�(�l��=��>#��֭�%#&:�kwL����=ȳ<��M�[��:��|2�LM�h$]=M��e�2e���q���n�FCn��p�%x6+��%�?����������N��q����I
���:�qK���ɚC�u��u+f���eQ��ņ���� xz��q��|l�C4���hhU(������f�xM�k����3˲�~���VV&BRĻ����@������h��'ǕNN�n�.蠡J;v�/p�Զ�/U>۴�������n�s�j��m[�o���v�ma�7���t�t@�����	�-{�n�59��h�OC*�'���[��b5���p?^x5��Ҿ �� <D��f�7�}�!-F�AnS�^hnc�E7n�]'O�5:�a{��Ģ��C��B�yd�W)���*>�1{�֒�6"�Y5W2���7��.	v��ᬰ~��9tqr#3��o*��}�h��J����9wV�5QMŚ����r �<k9���lP�:�+㭣s(ʑ�jP��'��m�D#����n/e!\,�8on��Ӿ������vź(�BY�'��!�?nj�GI�Dُ�No.���0=m�$�����_C��)��9��ߢ�0:fX��ع�1���=|��B���0^=�9��ﺡ W\`]��d�R�_�׹��.2��vB���	�
v�8)��P�".l�rߪAH�v�M�a����~\LB�
f�!�le50����q�g�A�+�gv���<������ܽ^�tÁ&�}E/�f6��6�q���,D�l~��֫��j�K���~l��n������w�����wPON����7$��H�"�Q J�|��U��L\[o���1/�/%�Y���#%W�4E&��r� r�C,����wq�`�_-����{�HٻV��zI�K'��\�OO���ߎ�%|ܬ���y�;�64"����U�u���d��DJp��($i�Ϣ����6S窧P�;E=
����>��������O�"
���>AA��]��436����?��2V��G�+x��v�~��WV�d�oV�|�9李Rkӵb�p�Ϛ��6������ᄘ��8۸'q�=����p���Cx8(e9)�ѩ1s��~��v�U�I��7��1��m�.�����`�\?��-��y(�+�7��Ѷߌ���cˁv��!���Taˉv����y�s&��b�	���
ɛ���w�#������bA��ۭ)��r�٧��{g�i�eS��_����|���G~=�}��iv�v2�>��x�1��Uy��o� -��nP,����0��8��X�W��S���z��,'�MG��=�����߾:o�o��?'Z=�-��,�1��y���mn�\�-WK�����<�Ǌ?x��޿O�M�B�b-��L�X#ԏ�~��dB������'���V��j�r$

��e6`#��t�V���ԾlW�]��I%�d_N|&g�Z�=t����l��ԉ��hp {t,}���(3zXw9��Q�Ϋ���>L�r�F�ɵ
�ß�RB�hr��Uto����3j�����AI���xVXPa�Ngwe���?��~/}��Ұ���g�!~`7a�D�|ᰩ?Uހ�bȞ�?�:��G*Fj"Ӫ�bw���,^�P����j�u&�v�)�@���#���ٽ�eI$�	��/|�.�z�9�h-��5��3rL�֔���g#������\����8:'܅,ө
���~.A�
��h��b�k�9����U{�tvo,��j�ؚrq5ǩI��;v�aDؗ^��Qw���z�����|�O��y�:LS�"7�)'�ԵԨ^>���B��წ{�נA����kK+���ީl*�[�Z2Mҽ�=��ӭɫ��Rh�d\�S>z��S�ff|���1d���V	y��rJ�>�����x�s_�Ʃ�����qz�m+�l�O��¿.��ON���4�K��b�v�ˑ�n���K�R�B�?S���������PX7������n3��sW�`]�dX����ӱ`h�R<j�`�O�����L���à��c.��y�q�g���&���H`c�}?X��%�_8J�o�;�0�@!�!��Z:��������I� �3�a>��+�O��W���+4��89wG�I�)*5�N�$]���� ���?�|S8cރ����8d/��j��9c	�yV/x(������^�`)���d6�bz�E�o�r�j�2���_��Q:k%\�����)ե��3�	��lv�~�A5�%���nH��v�V�����"mǵ&�&7�޹}j���e=LO0��͜��a\���/�p�LI��f^i�!�ഝ�R�pJ��
A�#�ֳv�n^��o4������y���=��.��"LM�G��G���>������H�:���i;}y��q���v��;�g�4�f�)���r�T��,�^��6˫$|\נ��l�q�#��ئWcP9���O��V3��z���Ǟ
m��wJ�,#��^2dHR!���0Y���&\�p�F�l��VW1�X%���4��=}���������3�s�������6�L$��M�{	7��<g��Y��c}���Z*�*����N����#-e�����n�Ǖ���Q����Z.Ps�\l@����'Xs����Z℟l.��� Q<���L��64�8H�q�n��~6��rS����Q1(���P��I�鯌f9R���m�yU���'ʒ�^�:��<��}�p��*�@��UF���_ ��O����|�:$�`����Θ�� �(\�Uw�9���AeMv��j�g~��)�
#v�S`)&�x�-`^�j�՞�h�,�d��Ԥ#�U2��Z7v}Qǅ>E��̷؞�X�V���i���WrH
^�#]"��8x@��������}2"L'�+m�%͊*�^d�H���r5ù�6�骜��5H�¿..e��7���hq�c�\����.�w�t��(2�k^Ť�/d;���DN�֊��"�hn��v?��׶�|�:m��:�f��9t��M�~(ƃ#��'��1!�b��7�E�l]��x������^��	�/z�i��,t���!c��y
|�'9��!���z{" m[Kc�{47�ɸ�I��U��~�B^�Y����I�~�\�)v�@]e�J�ꮃT<9U��X7B���MQ�ڙ9�N21p���/��7@p���4�u��JN�h��1|�~�ԪX�DO��x�N�A�T���l�-s~-�5�sH��T��\TќY${q��9E���E����#4�b)�P��N]KnIٮ��X�^�&��@k����g��ly�q��KYaHN}�}*$�Q�n����G�n�\u�`f)�K?�\�?:7��w�=����G3��KH�~�O�*�S�;��r���c@x��)J�jl���Jߡ������Н.Д��X�:�~�r`Zp��f�/��$D+��������CZ\��w��9Fr���ԽKش�?���KA��jq�RuFn��
-��]yn����'-3 i$����X�-$����e,,�Td��^�Ὧ�բg�2�K��`;�Zb�9��S����������YB�������$Q79wi[�^$��5��4�\�1+*���?b?��)E,ߥ%�S(��_bV��|�B[6�h�\���;�@;�ތSk/(Z���� Pݳc	$�n�T��+��A���N�s�MmKk��j,���F���A3�V悂����y]�7����g늦��Lv�ߚ��	��̍ԩ�@��\C����6x^.�m���b]:b-;|��Wb֪#Az��0P4����֫�vUp%6�y��Ҫo�d��Z����Ό񠳕A{���{ğmMֲًp�> *fs���]�?��ȓXC{=ҍO���ډ5�W/�\�-.���B�wڻt�����K-l���A|]]�1�R�4�Qf�`�����^�k�R;'�b�/Qg��B��P�y9}Ռ�U�8|��ƒ��!O���XN�mo:Z }ܶ�'��Xùhe=�]9���v��!��G�*Q~�/?1{��d5��^ߊ~-q.T��� ��v��^I%By�؉h��Ew���C���^��`�[��.;��
���Η"��2G�#�3w�����uK�� s6۱w�u��t{v߽�_Xɜw�����۫2�����tP"<]��/V7�� �����n`n)>�0Ƨ\�Zoq���G6{6P�Uc��0�H\u٩�+���6�p4BḠ���q����PG�����o}3���*#Hsߣ��ӖG�s~�E3^=q~�k�Kz�����0�ҘC[��ra��� rs^��-�H�o,c]�U�����Ƙn`�| Q 51�[��{H����Ko����
w���Z�+#[RX�C����1��uJ�;���Su����c;�^ 3�������8;�?\�{��\���δ�����Jf���eu���n�.QuG��D޶��˖��3®���a�{��ԾtL��J����
���z�_¯R���ӽqb����m��@�'�[��� j�_uE����-��B���l��;�5a1�$p���`ݻ��ȧ�dX
�4&g���_k������ظ3�z�d��w���j'd�"S8��a�f����Va��c֍R��������L�&��?�^�A��Q����u�}�p��-|�8fJ��?�<�̛�))"� ���P����v(í�zF1��v����h�w��j�{F�>�H<{odX0�*�����L�~zb�04�R��B�xs���2+~�C��ٸ�ٸڇF��\��'8�E�o���Gw���ץ#�L�bv���<���/�u&�\���B//��{#��Wk��N��U�H��Mb��ɨA����G~�/�4�!�U�W��3��Rz��̺訩3\;�t.����r�ry�t�N��!2WC��]�l�Z��a�n�jј�S n��Q��ݺ��~V�Uhs�Ĕ��F�I3v��X�~�nVu�(�_ F셄�I�������B�j�k��wgM�����:>o��W����'DdU��M�����S1jw�3�9-1;-�Mf{��8�v�cԪ�M�^�_��\Dg��D�a�!��+Dz! �c�L�Ѧ��Gmv�ᇠ�|��>+x�U	�?z���S�//ص\�׫��FIfS{=E�_�n���Xb�GG�N4�rka��uU>iE/[���A��9�z=!|d�8F�xd�n��9�9l���ۧ��]b/VPs�iӈ-!�ᱵ��kH���a�Β��.x�����
�N�x28j�VF�ב.ro�@7��������S�ը9�4F�?I<�zm�=�"ボ�g�H�5hN�d���m%�ݫ�p�	o<��sn���D1|O)�<��e.�K�$��o��/��C%��!M�	,��1����-��Y˹>�V����Ok�NO�E�4�䲂���(>�I,��ʧ$����E�_o~}��d_HT-��l$y�,:�;C#s��ҳM="�-1Fι'�ᷬ7�LW�!O����~���gƩ���l<39!��	�ڗ�Z�)�j_X���0&��z�,7��-i|>�ܓ`�ZL�ո�!�����5j��:+ZΘJYp]V��o�Jyx��1'�.f/�]�?|��Sy=r�K��-l����xZ䖭�v�^d�+(]]/m��tQW?P��;
��K�|��r��"=��GIp����q�W�'O]8.kX�.&���ewt�6�*$0Ю�w# � -���̾�� �k������<�� )�W�a��3�~:�3����-*ymo��:g0jz��k�4Z�g-�.Gzn[mU-i.k��Y�]n���W6Y����
	���O4~'RN�LW�� ���\�ǧ��"j��d(c��9*���PM:e��瀎y�߂C�U?�OSݳ9hA.�4��!_�1p��g�-"�܄baw���}-:s��i�Ml��E���Pʰ���~���qn�	�)���&����+y%F��ᄸW�'5bP�M�T��uyB\�����]����V��#4��9�YM�uhq�9�#8.��cȂ���&�g0?�_�*(�+[{{D�o�>�4I�\u#ĭ���SY��Gۙ��k�g�`���{P{?4�_�kq�bg~㋱���g�6���%��~ւtE���Ok��q/��9Tf�JBq�t�����τ�ѳ�,6����WjQ��.Z~�0R��r=��(F	����H�(c
��k4�幨K֣F��i��Tz S�4�__'��̂�������r�΂���(P\)��7�I23WpZ̾�_̤\�Yy�3�Δ�t���ف�+�.��w�b�H���t�q��7f�
�|��:5Q�%�y�z^<��`vd�%��� ���Jf��h�w��H_���>͓i�� ��e���8$�J?�f���H����R]ge�J�v�D��r�ύ`2��=Y���'\1���1 ,J��d�e�(VDTK���7�#��N�������)�[R/�nNh�sz�&k���w��j������A����>7<������a����*���\ˍ��o00&�)���_<u`��	�B��GO�pvOP/���JLgA!�p65����q��������%o+�>�{j�������PK   6��X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   6��X��D>  ?>  /   images/681693c6-5654-47c4-ac94-4786caa34b62.png?>���PNG

   IHDR   d   �   (�-F   	pHYs  ��  �����   tEXtSoftware www.inkscape.org��<  =�IDATx��}x�u�?3��ŢW�;ER%QT�:-Q�r��{�{lŶ�����;Q���ʲ;J,ٲ��%J�D�)���lߙy�3�X� � Rrx���3;3���Ϲ�����6Y�H���K��W�৯� �� M�m[�/���%���q�?�o\W�eeAܳw �n��-�Ć�����߄������x�=�]�q�N�<,|�
�ǎ^ܱ��H���P���ڃ�T��>�����R���`wW#㺤.���_�i�}^U���룿oD����?Z�C}1lk���4>�6���˱q� ��B'.^P�Ｅ^��?f�}�(j�eM9n{�	[[G��˪q��R�b{݁SʲqaM>��H��6 a����m�l.JJ'W/*�W���gj�ֶ(���Q�0zQ��T:GS��LbOw����͈���{����rܷߺ�߹��!�:2��܃=�yZ���,Ë�a������\���X+�m
��7�"����>�'���a���c�o�`4��ҧ&��2�no.�y]5�ws=��a���](Т��>��>75���o���\��է���������a��"L��B �[F��&�z��De�$�f`���\|��E��CMH�l��YA�r}:��Z|���jB�俄+CB�y!tE�1�?߱BQ�uK
q��-YC�5�i�]�.�h�U�|����P+H�_����&�;�� ?A���J�z�
|��fv��t6�ޟ�ׄ�$?�����������|��||c�Ɵ�=�5����|h4qW�*���6�qmF	���G���/ .綍��W��	!��en��6�]y;p]�>���<]����S��ѵ�������DU� ����s02�C��g-|���p˹e�������g!l~a�p����$��;+;q�M�CqYZ������Q��ޥ�]}
��l�[VUa�5�nx��!�m�{��p������0ޟ�7\}��}£�����ۼ�/����й�7�&\}ӧQ>o!ښw!��_H���~]8���y	oY^����,�� v�|?��6�߬w�+O���T�bx�9�t�z�u���EFP��O0��
�_������`+�]����	̫Y�ζ(|�5�Gె�����꺕���� ���W���/nT���#��G|f۲B��@"y�u�W_�Ҋ:un��uX��,�ۊ&}|B��ZKs��z��#�d[��f�ڷ�!te"�5�i�XTQ�kެ�)(����Ê֍��_M�[��ҳ.BE�bu��Ek�x�
,}��Z��F1,�uK?��P���7aϞ���GԨ i��{��4+/� �c ����ވ�ͿV N	2`�X�&,Yv��P�"З,=˷6a��P��h k.܀��buݚ��������t��f1��Den4<4�|<��e�sK�MJ8"ajB}�n��&Yjʄ}�lg�	yV<C2W��	ʳ|���,[�/�t�5���J]�-}
p�Ȩ�?v��K�L��H��5!�%!b*� �[0֧���aZT�p��g�}�w�)���F2���&�	d�4&���G۴ �Z�q��'��W����hܻ;ۇ��Z(Tm�T,��Q/'�b�3w��7��Ϗ][6b[�Vc!*B:bb}JV�~���pɵ�����a�y���a�XoGGLl�Va��G�W�QQj�����҅��:4y>��H��X��=�̔pf>vo} ���q�,KK�t�#�Jl
���;�K�Gx�OD����y����i�}�ī�Y��� 
6�Vqdk�v�j<��[�%8��/z%�����)�K^��8�AA��2�%��,y`$ea$n���[/%�+q��Pd<�6�%7`��ÿ�X���d�ȽG���|$;Dw�w7(E����(��"�����&���k�Ϣעg�,<p"����ǖ��V�����}Q���`�Ǹ�^A��:�B<��]f�ym5޲���	���[î~�fbj>�_�,'�N��н��El=����w"f��OEW���y�R����M�g�Z4���[^B����Rע9Y��^=�?�_x����FF���o'W�$/��ɸ~��C��,��|�)|�YQ�w�c���w_�I�u¼)D� �b��-�1,H��#-b�/��n�}m�I�\e��
����S1-��b���w�+���؛�J~GL�[]�O]T����_��_�\�7E,�K�"GP����u���	�*���u���O����5x�X��P�Y'\��w,�Ϸ�� G�/�Y���_F�F��Tb*,}�uy�xy5n���]<���*|��P�f1Ɠ"�Đ���ը-��C�k��lӻq��A�JhWq�޾���bp������B1�I��s?|�B\/�m8�(+[�U���v1��"f1mn��o�P�va�4��u�ů 2����J) ��-E�x|uѢ����}Gā��֍G��7/ă�D���|4������GZ���m��lX��pRܱ�/�'���R������o߿D8t�O��hRN�m=��1d�C��>�����m6cT�r�b��Ou�5�h�i
��kg/~(�mȟ=2�F��P�`,%�u�~w���qyM9M���A��K���k�*/�Q�~�S�hPy��x]����hJ]IXʳ'G�	�}
!�A���^�����I��}���#quۏ�u���!E�v�u��I�>�%p3�����q�Kyݾ�(>p�a�����$�bB ��t�1-���e�Fz��!�y���`�PSf��߼�|C-���^�����Lѧ6�gO$��p��g��rC� ��>Ǯ#a��)���<���I8�"=��S�C++��.۟��Ag1�l�<|��u�'a1C�Oڦ��3mn����Z!TJI�	�Ol41����&k�i�7�"�27�sK�	�ØM��o&����/�;��9n
!I[Ǌ�!|��&�-��@���0O2C��M����芕�P��h6�q��;ѧ>����o
ꎃG�9���>�rs���4)�N� 	�\��W'ě�g�6�R�ki���k��I<�>��ӌ��ަ�(N�l��(,Y
� ���JA�S��?��]�M	��u`�у�f9V}�nV�b�(�K�c���O-��<�Z����Tr1��7���u��4�P?�s�1fF�4��V�P]~nB99j�9�"�D\�4�g�jB���p�h�|�BL_/�z?L1<�i�>�!31� �TH}ک^��Q����S>h2';'�?��L���RB�<3�^|6M!��-�G�w��<�'0�8Y]�|�DW�1Rם�&V����|�Zl�1�r�E�"�r��O�Y?��/�)��O>s�
rst�KnAϊ����969c^��]��(ׇ��a��\}�C��
!\n����H�}�twU.�&�\�^C;�<"@��F��"����tw�'sޱ�#N��g.9�f��@�f�����!������̜T݇���c"K��D�1n��y�5�$��i�N�Q;��=�S��^I�R(��Wˮ�4��J��u�=Iy�֗��M87E���644�Dr)#'cٵq�:��4�"���7d���K�:��2�! 9I�h�̈́�x�_���>+��r�ײD,������Y&S>W�O�Vݸ¿���*������9�"�%�){*���x�g@��Y��/��c��wc�]���H&x�;ߊ��K���� �^W��'k{q�]w�A��/++ŵ��>�9���5c'��p�9/R@%�n�0������s�0����AH�7.���?�H$� LĿ�������@_��=����J�Al��B���X]Bii	��[P�O O�*WK�di!P9��Dm���E\͛��d?a; ��,6�#�IB!8i�K��;��'Ї�s�g6<����E��]
��s�X*��v�8���\|��O�8h`0Ǔ[��x�I�\�
����^���$�`$U��@}�J���̿��yf��L��4���k����-7Ll|������h�r]<1RRf*�%C�`�I,��c��DLh��-�����iCi�����[<�қ1�v}����n��⊍ruOo_�o��$#z�D��'%��]V� b��!>)*�� Em� ���Y���1T�ּ1}�eSLL��1�}��]�cV�fFyY��5*V�Z��#��(��8,��!�J;P��t�ir�7�?	��.��".bӢ�5>)(�[�<7�坐C<��	A/X>��"�|�䖧2f�Ī�Y������2���C���˗�I5�e�I�,���>��#ibT�S6f�\�S��0��(�8��z��N��23m����K�8S�*�R�H�$(��d�>$������"�D��V�Àf�H����s�z�ODD�^�-P�)'l�G���R`pUy)"9�hL�)�ז5�ׇq�����P0�E�cǠ������&�p�,�nj*�8{b���ߜ�^�#� ���ڢj�n���◝�t	�Gr0��f)c~�@���}~3^���8f�����T\�zi�>�{�,+Kt�I�Q�������\�b�����񛿄����x0�=X�>�*�G�>�E!���Q��ڑ4�D))$�� ��ea|��w"�`������Ư��ʰo�L|O�?�����9C��@;�'����.�}Ǆ���b~]bb�����N&�J��ʠ[��!~���A�rJV��1���B�WU�$FOw�*�p�D��.'�ru�v~���G�1|��a�~d+�Ǭ,z�@��á*�~�|I����q�?�6���gPG�U�����)*).�֣�%3$�L�_���2�T�oSot!��B3�O�������Z�"ĺ�
9��
�D��c�L?%C���P��ʪą@��Y�ɢ�BS�_��d��sޜ���A�pL��1G��r����Ю��;�E(h�az�3�l�)�����$g ��j�V:Ru�<!2�/{c6�z��%���?��0D�O�~����$���4r�B�AX�Ō���+͘p��N�����a�ј9M�n1%�Z��a�f����b�-�5`�Y�v� ;�5a�l�oj {�?�H���9^������sވx���8v|P����Б�*��/~�Z��!;2]�P�$�I�� J������?��ؙ�"�!�8��ԩ�h��˜����b�מ2�=��Ԧ����̞d���B9/��D8��?֯_�b�!ñ6��5����� FlACc���L�k�C{�Y��p4h^��̇���'�N�,����.cbIk�U*�G�`^n���m&�A���ƺ^9�'�<[S�V��D6��>P3�{�W-���@ ��������B��v���9�^z�c�D
�ΰ�qg�o�ch�� ����	(?dCQ=���xC�B̻��S��yQ��2-��jq}�����"8��RN,'9��{tM���oR'�Q�P��a4Z%X.��^����kUb�ރb�3ڕa����#�eH�8'��9�B6Mž:�W��+zȱ:�C�DpU�[�@�����VN��m|m�h:�'�Чh���d�=��c�4��v��$�M9�h�Zu���\�Ԉ��/��M�b��S�Q��pj�5�R�Q/T�/��ADcLr� �T�6L��'SɄ_y���3��t�$�]i�PGܳoV��u7�W�s�38��rǮ�������}�oN��C�·6w��Zx���l���zm�pF���D���>q�"f=��\<l.��<�I��s�|�p��X�<��ʩ���4���F$D�)+����,�O����1�Hg� �χ=�Pk��Β	z-���M��訍_�T���:�e?�]I���x#@�S����6��g�JS���N��G���H�8Q�=a�n�������"�����m:���t˩5�(i�`��b�%!�X���Z`~�K=�ŵ���k��R�5�b�7����F {~É>}�gڔg�=#�K��&�I�H����BW���ocK��2a2%�8�0TpAA߸��ԕ+��VC� ��y����tI��n��m�c��z��n��*�H庖�Ѣ�]A�_�|��+?����=��+)�,#��ǅ�ˌ8�����cݝ_6�)l�Ϳ9����n������:���@�>)�s�8��`4�k� ����'B
w���R_�aw����2|z^����ӥ�i�p_�kꃂ�E��K�j�Εa��� ,��U����w��]��PQQ�?�)|�8�������Q����-�s����yJ���m�����&��\K$�tA�%�㐑n� >r�"�d�&50�YV]GU-�.�NUO,�,�5P�V,LS�X�GI.�B#$JC>Ya��ExA=����˔:�A?�+K����8��b5�ŕ���>~�1�.fm�p4�$��&��b�gOmc$iT��MmL=�/:�}�#2��	�'BGR��WL~�`�D�<V�|;<$@�ca�9GC1��;��:���z��dO"+>����=τ��^�F�Z����>��;�o�o�0�O��������v�����&��w�����D�ﮰ�SÝ�\����Z_$�O�߄��Ѵ����΃�zƠ�ht8z�-��;�9�vv������X\��/��	��϶��av|���l�q���;�Z��pT�S3H��Q��4Co�v�s�4��}����Ǖ��/����a�M�'�$�)=�$~(X%��hW{�a�)od ���\����ҏp��c�n:!^��Z��s*u�hg�0���-�&b���qaNu��9�\��
�{���Ԇ�i3k�ge���j<�,z
�?�RW��y�*Kh��j��A�����8�-�o*y�,�����\R��s�)d���ˢ
��֧~|C�
��3��XW$�����Y	���7���}��(
jxZ8�p�`��Ѥ�m��V���Z������+D���b��AΞK}���ۈ$m������f�����5����)�����j/
īX-�a4aco���i�Q�4��*�q��H��"b�K>��L��yȑAK))C�b��2�~�s������d ~�=tRq�{4��S�M41�n2O%��{�L��&�s�EE:�_�����E��g	#���L�	�.$qϵaC�!pk��6����zC=|(ncG��t���R��s��X���y�e�AQrHwvD�v�X�q���ɅE�mn���s����AT��{��ykX;�=�gy���s��cخ
j4T�bs���H/�O�]�(��2]Z��&��Ԍ��-:���	Ǻ"R�%D�&�!�/�)�gT ��!����&��z�==��=`_�D�ʪr�YGGt��q8	81�����7�wb}e�e�Z�h�B��	|���?��%U��/Oq��rϕI���-)4�^-DMvOJ�ab��a|�r���C��j-Q���E�g�m*����/��a�r����]A}��HSz��A���(\A��ȡ�!�A���}x�1��;��P""O��C��8�T��.�=�!���,�(s8e�tB��O0�rv��L��?���m���u7�W�De�t����~+��� ���:�Ƣy�1�i��=���z��8U�v�ݏ�<��o[�J���P���w⎧~���G�kQt�`yr�����PW�T'��Y`D�3�2A�N�Q<]\#��d��VS��Ǵb���m�	�u��y��*!��4���U�w��8r�D������h��9 s�l/|G�O��ǯ	�>�K��2�x�m�{2�E�I��w��&XPU��V�1'j^���M�5u�C�t�vFhJ���7��v�O�V=�B��WҎ	PfWH=Uʋ�pѰ��
Ȫ�E��!�4�ISe:��@�ꛓi:���8��@ �J_�	�����g3�v��椒2�<��we�݉c���ZR��[e��jqi
�@wa��h
�)��$w�j���Y�s�C@o�J��J��r�;�˰4�:s�rm�ǚ���4l��N����UY^.�k�����\g��)�U_A~��,Q\���҈��	`ѢE�$�R���=�d���k�z��\�%�O`�h��Ԝm;<��mV7��� ��v�U���ը^yeV[Jq]qI).���*,�1��9&T���q�57�yN��mC0;R����I��g��R���q��KǛF`��QYQ]�7��3J����"Y�����#l�<Vxм���Nۮ�d��w$���BZ�/]D�?I_����z�櫉�N���'��}X��G[=17�I�kb���Q�%�4c�]�m���e���H����h���6�=����f�r�U�or�{�e�!1��Cfڴc�L�[��Ox�v��NQ��SiDؙǎQsf#�S��:c:x����{�������:ӎߴ����9Ӳo�:$�!�BNe��DV:�z�C�����0�������v<�׳�� �7o��t��K3� �4�t+C�x�"��Xy#5o�|6��,�{��O�R��Jr4�.�Fj�AM-����A
�ׁ�K*cJ�znL!������m���v��F-�<{�aym<�80�N���eN�=�[���"�By��z=��ziF\�~��ě�j�/3j&�YNM�xJ�O�RW���:��L����U�kX/�G�^WU���r�d"�y�Id����c�Z;���2�
?�}p��9HL�p�'���:��Wj�^��\7��d2 �5����
a�SEH�%BXL��k�f"��D��T�DdqAhe��2+�I�Mgc�y�R΂?�yU��i��^�3D�v8	m���b�H$	�CnZ�S����'�%* ڸ���!��T,*�r�T�~�F!��)Lv9�t��\Q<�LW��ϴ���^<j�A ESxhR�\0��e����1S��~����9A��V.���uRr��iX)�&u1�Z#��)�p�ٹƴ�NE�24�u��
'͓ ��+��3�:l���C�O��y�7ݖ�D=qs&�8AV]Ѳ"Փh��/�F��I�-(d*��-m&��8��:��I����<��"���d��\q�g��,���<�$saKqs�Y�A�BΟ.�d&���{�d?&�J!k��,zL�1�\�a2�i�J#h����N�ua�m��=�Q�ٽ��r�7�Rp��A��>M���Q[���ݖ���_f*�t�S1-{�L�!i+��}V���
�i��1WO�Xw��&3I�\���1����.�ud3�uo���/�m����P4DW����XK��4ԫ��#�c�<�)N1�R�.����O��%<O�we��Rf9'"���0`)r:\�L�L2A���U7К��eG��
�暽�r᠝2qN���ɱ�������EL���x@5-[�ɯ,b����|r��7y���t�a ��}1������9f�3�s� �O���1i��Ǐ�\g�RB�E""��L.f�,Eke���=�#d2�Ho�鞛]�%_ �AJ�gˁR��"�R��ĸT�+�h�Pw<�2fyёd�Q�3���9�x~*�|
q���!S�n��CrsI���|?j��s��-,}��H#�Ф����� �>5���Q�B������wY�D�E��1j��wf�OD�bXs�*q僢6:R��E�W��4ʤ����g�L)>�V��ZG�QD��
�"A+����U[R�Mބ89����VV�q�B�v��J�SD߇���ŮO��6
�P�6;ʛ\q�<��t	q� � ǩ k��^Z����Ŗ6Ag&[{m�b�^8)���b��$b��sj)<qV)ȣb}�)��g��ٮ�B3�I��q� 㒺|����Q��:���2��L�,ۇꯡ$���c]MH]�rۨ�~0�J0S�J�����E�>�����1��j("�;b	W��s�{8+4���2EU���U���"@�}8���G�cǬu�*�E�-����e�N���>����/���<��g���PL鄩^�̳�o�dTXb��"\P��A�+��5˅�m�{ЍSqL4.X����� �PLq�Dȁ~��(�V.D�8����4�dr�\9��k6E:��I��$����3:Y:�ku�1G�QܱP�ѕѼ߯�JL�=X<d�;�1oymO$�g�Fpò"��g��$�6R�cx2z��M�)��@�&�Ϸ?@�k+D���5J�X� ,��Enp�	���B��R4E���Gt����58��XC��:Ǵ�X'���%y�8���ܱ�<U��Z��#:�}����犕��쿂1v��Ek�i�$n�D�D�p޿�&g�n���~��Jr��^���:z%A]�G�� � V(���K[H|Ur/7�<ѫ
'[��R�^0+�8p��#I�5/J"[�D^��p�]1$e�3F\����(8I�?�\�TL["��Έ�X������e�6�]�OR2p���P�:{[��}=1�U�g�`wWT=/��*"l�CQ�#q4Ct�Kh<��h�Šj	Y�ϗL���3��tp1�Ef�Cl��ܫ;䱪���ci,z���q��<YߡJ�/�m���|"Ǔb�%UM][��Ӎ#h�J�Y�)�V��:�7-�QKq�J���yb�qs�R��M���GY�ٔ��c�1Mn�G�K��s�:A�˩Nv�ɹp��i'�-�g�K1n�5�t8�w<� U��[��c8�W@J��Mм�v�SH���j�yi���\�E%9��$���Y)�O����)�2JP��y�_WN)�+.jq��Q+�a���HH<Jlڎ� ��ߦ�ټz��"f"-sm}֭,O�yΜ'F�u�rNF�Gs�Sn�#c}��ջv�N��bAE�"�"�V��wμ\<rh�Ą70�N�4u��+aE��%��<���ǡ�r�t�`�c�q�Ǘ�f��w���1|'���D�S�b�]id6��F�t"n(�#C)��y��� @����pS��G06���Ή���r�RǱ+���*�Is�C�T�O�ҁC�5|良���F�QSq�����Ն�^���S4�t4��*�	���s����Y�D���W-�w-&o���-6ƊZMkl�����|��hV�~<�C�M�M����M�N��U�&��QtȜ'Z<4�� Ԩgt��ꍕ"��^T��Z:y�-�6�q� �k�S�Җ��/�?+�v�����c�+��p��
X�9�#ӛ�$�g���Z��>v��p��L�s�T�(���o;'*H��4�nB_$���vx̤��(3��C�|M<�8���]+K�v�]by	lDFe�S�~�x弿Wt����;�MX�d�KZw|��e�'�C�&$0��<�7D𞨋 �E�(df��v�5.Ff]d9�P���1������Ds���C��&r)����V8 r6���WWW�b��Q��("��N|���V��B�3�!aE���	���(���(?�A�p�T�X����A @�p��*V�9�D9�9v����0.��shg=�΁r�� ��"�����NiN�3P<2�8��F��GM�!#r��I稩�2w���[oI "��=s��t��c���\���}'R�3�$Rw�����m�=�L�{#�#gcl��ɋ�1ǌ�K�\�&�$��r�5�?{¹9Q�CU�ND�"����8�$��㤽X���}W�s�5Ǝ����8�t��\%��;oS�P��ꓙ&��t�Cd�W�CI3�������&',+uV)��ȭܧ�;�,�$�ވ���c������6#�3M"�'|�ͪBQD�S,1Q�S&wV�Oq�Di/+�9bI��Z^�Sg� �g�jWT�F��)�B�K�T��y�������CD�sD����S!:���/�]����䲑2y��L'j0��r���L��sH��5a=���F��R�e���
*>�q!RS��/#���\�8A���f� �d.1y���u
��{Z��@�&Q
����?���1���*��v6|�)�c��9&9."���=�\��B�k]N���:?C��U_� �+�l���I��r�B���6��f��=��1��+��@�CS�������K\�Y]�E('�ͭS�[�S��Nl�8�H��!��g)T��4��A6�r^�M��8�U>g�a��T�;�˼�C4LΣ���.�r��Tnju�u^Vb��4ƨV��.�A���d�$8�x:-ST͹�N����bל$����b����F7�cE��|�Ikݼ�����&��B�l��+�^��L���$ }�T�л��^���:���"�吺ʔ���R������F�)�8c:,�צ3��I.��M"Ӧ�>':���&��?8�^���cҮ�Xu(�ܱ��@����M��Kk<��&�����2g��U���c8�\A_�B�gd7�r�/�|U�J`�j��r�CYk�:SN@��e���#��*���?a�uF�p>�r��Nv�N�2B<�Ek�J��f{��}*�J.!�Ѽe:�ܦ��2������S%�9�'�E/|Py�cps�|S@�g��	gb�WnL�e�0I��Q��4�i}����;t`��ϝF��Dz'�s*�8Y�WS,Ѭ���p�J�kEC�q3anɤ^CNbZN8�}����309����>�:��aV̳-f�f�	uE���I��.��gPQ5Itq�YGIg��M\�$��A$ЙM�M�_uu?/�6x]�+"f �5ӵ���Q�p�W���!�7��ʞDD�q�%	��8�p����� f�1%�2�43�D@.Qi�}Nu��NG9��Fky&�wv;��J�ce�i��ƴ��P~C-3�d��Y�}b'����l�>17�M�>��P-*/�}���Y��X*	U�C�a�+�G�cU���4���ݦ0��!lTv���(���'�K*���=��R>��X6���袧�T[*��Y���)3A�X��)\1d?,�a��^��,�w���0��^'���E{�#n�ZAE+�����>�vJ8�����z�7WP&S�Ӿ��R<��R_��Ϥk��<��&�TYt�Y��e���z�}�F���ey���	���5ϫ�`}��7=dL��P֩�t'2�P���0}��44ϫ��01c�1񙓝;mY'T�odx͋<�֐���)E�	^��!�v�~�e4�xf����i'nSI���!L�qvR���ʛټ��:�d�g6�}&����x/�"�N2����X��
u�N3�b�ݎ��fI�;nF��+����Dj�Y�S�c+}(W��c�Z�����,�3�����}�U���ѱ5Ь�e�����5�ډ�2KR
����I��5�:�(���LΒ��o�p0�`��NOXR�B�'�SX�o�4��Q��O��y�:�vS�B 3����ދ?�x޵�De�on�Ç�������O��޹X�>�\G���mNb�'�"�/+�W�עs$�����ZT)�?o��Ҳ�Ԏ�~��w�g�Bl�x��y�o^\��\2O!���_��>��o_Y�����ُ;^�QH���$�s�>�G�I��8�R�~�6B�^���ksp��R�r�%TV�7v�Л��w��%�[76�,�x�|�jg
�;n�܉��է�qY�Ƥ6����m�~��* ���*͔!g1�+O��޳T��
��C�L�#gy�/���ۨ�~�X.|�a�)��������}N�$s����� Mu�y'�h�y�K�:��7.��I12�0�\���o�Kp��K���o�FQVЄ[����_��ԃ821W�f�%��"4�Ǖ(��<�L��܅���Fݟ���n��m����D���W�êP���?~�"l�?��)J�)�8^O1ű'��B��_j힥����e(�ĥ�������W����w��l�,��w/���.�'M�՟��^��:���&���&6���P�߾P%��գ�0M'�����
��=�*�g"H��xa25S|X�I@���RE��3G���U9���mQ|Pg}�6����G��j]���S"2���"�&��Ay��/���:9��Ib&�Q���j22�g�7E�p̔Ɓ;�+uK���E�E��t?։{��s��~r\���M�6��x�[��M6��>�)���1��<�>Ӏn ޻o@�R��EG|�:T�����l[%Y?xpI��E?�j��������{Dq
E$�p�菜I�����JI����|*U�D�l"7�B,�o�������v��J�_�����_�E"�9A*рOOo���VP(��T�g����bi����)*�+b�Q��XS�RN?x^9^hUȾ�*{Y��cD7�N���~,���xE5��X���#��gu)>q_�B�gO����`O���l��c%	cgg����-dr�����d�"�ơ㚊�"�8R�CB���I�)��N����$���[*q��P���*��xn8n�<,CD���W��[�T	�o߿L=����̯����O=� �C��j��G���fU�N��ߥO*�|�Emh3Q9���g���˰�����7ԙ5��
���dm�/k��]W��U9�9_�����F�F�����c׿{�MM���\��nb�g^2��_D!�}��Fu�5,#�=�0g��±�:�~�_	 Y���OE]��ͬS'`���#J�(ȉ�W��LGr�i�K���i�q9	ݓ)c��o��5�
���lD֗oU�3ǭ!a�0ӎ���"ޓ<wR�x�2{�a�����٦���?<ێ��ܲ��W�s{�hVb�xm���i��3�9oOs�#uzf�T��[�55�K۸�6�w�"��$m��xjl2]sj\��M֜=SRx�V����Y4�wwG������h�09&r�L��3��YZY^9W���NS�M2Փ����~�w ��7�(<�&�Қ�\�����@��>�s�)K��[�����3ճ&S��-�p�3J��B�D�h�T�P�y�D�ԍ�v�J$�|a^1���W�+�T�����Ɯ)n�}������39#cR��BF>O���@1!-���֜����[3aA�e�)��_81��Q�b� 3z�hl>�i}p���v:B2ݓY�\�$���`��?��+sN*.a�6��^��8A���`v$�Z.�ᆚNQ,� Yv�=!��gU�T���d0&@3��Y����u���@�b���EB��Y������k6kcXf�d�;,%�X��0`N�C&�q77�2c�Il����l{�)VÊ2Mm��}9xn��F�6�-F��,�c�1�2��B��$h�{�Ddn*L�9U��L��@˄+����\��ؘ��N���f�EW��8N��`:-+"����SK��}Y���49x*y��!p	�P+�R�������csӎ���-�BB92�Y��Nuc����2�c��0�6�����lSz�[�MA�yZ(�cL�Ζ��z�Ck��&�0M�������i�\��������2��\    IEND�B`�PK   6��X���&  �&  /   images/6cd43c8a-9a35-40bc-b660-85b087cb5f0d.png�&wىPNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  &IDATx��]|T����]��{B� 		!�"� �X�wł�{G�Y v�+���� ������4�JBz�����̻;R�@�?�����������ݝ��=)BA��D��б�q��n�b6���2�jU?�h�8�n	b7�C�ig!p�(xv���My9���g�����h��p�DQ`��~��6�ix��h֡���`��Dִ�Q�b	�z��qQ�^Ј vQ1�<��'��Wlw�z�#x�ߜ�^���ǡ}�ES�]�"1_k��@��%��q�b��H�ht:��F��N�:J�v�ZDw��F:�����q��>�}t�Y�;��y�]���Y|/�􈃌��	1�V�>��kM�~$Y�{�$B�W�m))��0���<��*��0��K�i�O�~2�ڔm�V����{y�;!	��*��s���WL��1Ki1a� ������a))j|��C����x$Įs2��8�Q��DUЩg«[\��}�o���qp	?؋��˕B(���{&ލ��'#��q����Ly�H��*���("�M��d�R�u�w�݄���C͖��z�Ytݍ�n��y�t�T"���A:�����ա�Ko�Z^��)��$�qY4+4�&܁�Q�#��˙> �-J��v�p��""a..�1��^Ux�C~�-�zA�o�
��Λ�F�$��Q�oE��!��9��;d�2��.���a�J��1�
��܁�i���	�ݹ]�:�!ѫ{<Y|1t�py
#����g"���P��o�}���S��K�"K1��.\�ӻ/��P����9F��}ąv�A��NV�(_�U����
�?��K?�eh}}�C)������Q� ,C�E�oc9�Q_�q�x�>�z�h����CSU!b�^[��A'�>s���K����	�g;���\\[m!�TxFǒX��f��'����>A��5�5:_?zF⧼��%_a��z��}�.��+�!���P��;қ�Bh�C���{(]�	/��]�߂��[]��p�ՁGp�&�}x��^���_%Q�Klckƍ��Q]y���93� ���z�Z��?SqjEę���1�oi6�l�G�����t��/�����[�Cܤ��,�VtB�o���{��Mt�aQ������.:�4A����w�x��AT�ɇp `���q����G ��Y.ǛA�!4[M�ه�P���h��p�.}�c(Y��π��P����g�p5�nB�=���� ��݅޳�ӌ_����P�F��*�"H����P&���^��1��!�%�QK�1���Kڜ������ u�D�9��
~J"�v��U<2�ocW���>s�ZU%�3�Y�:9�É<�eW�pH�n�\���(Y�].�=�|;��HE��R��(^�}�-!�T+��l�Ju��uD2���u��}J{�s�g�W��_0v?|�)���x|{!����I�3{��X&�7늲�V"�	���vx�8,�~%DT ��{��Hg���㩩�L&Cșc�A�C�O?P�4x��٦s���xV��r�z��|i��ؽ��K��VN�]�E��V�"�T�l��[�����f�1;��	�do��|���?~��6f���q��P��IE}�A��I��ɽ�������<+������7j�B��WA]�zNZ#1rH!1��'E\�~�6��M�&`��j��U���c����� �܇�6r�,X��G��RY��?U$S�(M�=.�U��L���o��h����W�$�����f��� %+��s���n�"���W�V�i��Z�`.*�	��^�q��`B�Dcc�!�Wy�����R~�~��@�3BK��|y
z���V=7���>n�����j�6��TF��Ev� ���Q?"��f"PSO\&B�۸�/�qw������nӟ8��5������J�56BH�̷%ҍ�7�w�,�5�9"�r�s -�4�͞��-�;�1oU��J�D���g��ǐ	8Z�~��.��X+���օ�5/���+��%d��E�#ޤ��$��=P��+��)�9�;��fs7���m›��hVz^/&���I��hi1����2:�lb7�=;d,���Oΐ����M�Ë-��"=7s�H��"z���7"J^�a���[��ތ`�	�Ie�gsX�l1
1����ڋe��	��6א%�=��&�YG6y���CaO.�;Y'�a;���k��eZጢ�dd�<F�g�D�e��u�V��Q��F�:<�́;|�im�1���w��=��TC�pO�d��֢��f_?4�Y��*z�[�:��U�Tk����M�a���,޾t-�<x��x�eי�X��ϝ����C��ݪ����f�FQ؆&m�fm��9@[g ^I-��S|6��׷z�t�������V �NĹ�����!��@3�Z�5M�ȧ��C����6���!$Z�X�l @q/���&�2�Wm|8�
G� �(o�r+6�M>��~�8Q�2ω@d��[�u����(鑈���+��	�����u�i�a�:n�������z�0b��cWNOm:jc���5�;����$昀V�'�A�Vx>���kuB"�ZXȒc?vU���&"��o����R��������;�!a��m�b��Lh��c�[w�˳��o�#�s-j��@}F��������[#mu�3P[�TD��l��܇���S��eK�y��Te�b�#�(y��{����\�Φ]�V�4EQ���]�r�v�!��\r�A<yFgf�^�E��Z��/�&7���0Bm%�����r�6uJk*k�)Kq=�g���?L��J��*t��b"�ǃř����kc��$L.�Lӹ������:��8A:�g����E9�|�f� ��V�p���׎cD5��B���n���7a���V�#����� |��x�u��Z�k-��ʋO]�������Mu�������V{�a�����ڕQ��6
:K��x�zD��zD�$�<Ǻ��k=�u�l�?�:�P��b0���Q��o�|���<L|���R�D������"P���Zq4@6��=~-���IkǠX�x��ެo%��B�o�>����j!�]��U�i������6-��lda5���Q�����뜑����򬩆We��fE%������4A�VXuLV_���f����R��8:�9�	�����I��<lH�I �˝��8�o-�=��	}���I%ao�YG��ϑ	���q��*r[kr0�5�]>�O���Ǒe������I�L7y�5-/t��6�t��͑��AZ& sM�x��ax���o�-Z�G4GakQ�D��ec�`߿oJl���#�j��too[�غ:��XBF�/��&k����~�N�sNg1A__�����w��jr�u5�6��'��>*�ə�v9k6�>8)T��Jׄ��ގ![3�x�q�N]��y�(� �<2e~Z%b��<
���
RygGߕ_�2/;t���c��3�����3�9vT��g_&;K8�0��y0�Tɞ�cw�E�X/�I����wl�4�t�r�:Q䳞�(�����R�'���Ɓ<��^��y+j�$�YoЫajg˱ѧ�m*m4"[�rC�ƽGVhPt"F��n�&�8�P�v��Ѧ(�>����6�T�|��y�5M�	��������<���x��Q�Ǹo=t��g"��s���q�-�-�z>���iO�(|5>ch��9��:�a�# ��fg;D�����Q{B��m�n���QϤ7ls)����9�N�ڠq�v,C���,�KR�/�m�Nj�s�|�5jc�B�[����E���u����Ӫ�(��X�_ ����������p�ص:�l�C;^������U��e�6Yf����o�\/m��f��7`�6''0Q|�K��ۅ�	�Dpf�X:��nk��E�}'BD�nsqBSKOU��K���-8{�d<P�G�m�|��\�g����GL���$z�%Vu����l��N�����{g���dp� �����q�t2�\�C�M�x��A�!����$����9�&��:A8�j�G'#��%Ki��P�e�9�����y���V5�����s*��Dg�ι�^/�1�Q�p�$���?]o��O��ZU��7^B��EnsLq�W�f��:??�r�Q�7UM�vrV�@�X�S=����7`02^xZ�݊�W��g
u3۹�1'���$��/��Їu�
����>	����9���CMK�i�����&9֐�<Q��d��G�Lᮭ�� RfA�÷Ot��Z���X$|>[��*bG�9[ �;�Yv:�����}����a�}�����\��R
r�����9/��]݃'�z�C��^.ig5G!Ig���I=$��d�p0PS�"��+�'��m���E��Ks������������J�X5�w� %,�>CONѠ�����I69�2���$�����	�����"�]���[4���z{K�����gLw(��hI�_�"I3[/o���q���u���C��$��3��ax2toL�;Hu�;��|���C+b��K�F�cF:��}�������[Kf(�պ F)����
����C~��RQ�����s�U��� l�E��-��'�w\�fcc��l�3$�	G����]��h���?��
s��	arP�ݙ�	�yy��n��O$�����N�|��vۖf�/X<�<ѷߧ�4��镌����#��ǜ#"ѻg/胂����ٺɽ���SwH5���ԯ�u��h8.�iݗ��x�mߞ�z���PbU�r����@�!D�")N�6�%Y��[8q}��/`�uK�F���f�� �*|h�������ۚỎ\ǃϜ�#��e��3�eD��f�4�Q�����`�G:ɳs)���>bx��s�_��~���jW?'�� �@&h�h���Rja�c��
n5�턈���>}����!*Z�%Ί��̤��8���O8	Q�ߢ��͒�9웤O~T��p���^y�'�]�bT�y������Òƻi9�Rg7[T������6�{F�L�y3�Kn��$���mM��LǮ��)/#�a)/U�2�v�w�d�n:Ywxu�C�E��Rz�o����/�J��jT��S3뇑�O����_�x[uI�̑�֊�f\�-�l�${fN=�BIz�U��b�\��8��N8Y�)q�2�hm����	���һok-+uzQ��F�<e��O6����w"bx\��f}h�_t�p;{�� )w�u�X�T��c�=$Ҙ�\ˊ����	�|�H����������$��8W=W�a�/��Уu��?0E�S���҇�I����Q�y#l�����;�-��.���m�b�P�r�T8c�P��b\)G��s~�� 3�p6�}���U��l�"���p���o����<�c#�s����_��3�M��-'���=�Ԓz��y�WI�p�/�܋�k�L"x1J�|��O?��q8���Y�:�5�?���fI,�ݞv%�f_�O#��w�G0���Ÿr�]�B6�Ѝ*~]��{&�D;O ��D1 ҟ�=���A�ƈU�r:�;$�:�I{�A�:���r2���L�|��Z�穩��� ),Ɠ@ә	��:v����%��yYM�|-�v?rbɓ;�2X++�;�-�cܕj��XWp�����f#}����s�bkm=C�/p� o���jjX6贳ЅLx�p��K���
>��om� 4����rA\��T����Ȩٶ�U1�ЋV���H�pҷ� ��X�'�gS����#���M�;��<��b:��â��n>��w�!᥷�����#��f��Fc�<�d�q�M��>��ﾕ�b�uv�1,N$�4�S��Ƣ$�g0A�ۯ"��W��^ATD�|�HLY�^���Q�={�O��f�(�hH,r��g���/Cכ�S;�^��t�r��=OG`����~�|�;�$]�O�7o?%4w�R.�#Q�o�R����}ơ��z�#�G�>�A�ѷ�t�ٹ����H�'�=[�~��x��<C^�a�Y� �눻R��t�y�n�R1�FR�K�� !�+�ɠh������}di]�H���ٍ��Z^>��H�q�|��?�C��_����}�Q\��Z]��K�����RS7�̱H��RW-���t.n|�jA�.���2��W��=�nKE�����׼[|'���WjUg�c=�hl�1]��p\w�k�2"ي�q�<wgH�;8�^�.4V�`�p�\u���n5��or?�����u'�dr�U���N�H6v���1�.;o�F|�A��,�hӺՇN>�E��}.)��]ĕ�KH�k�Ӽ}+t��6m@��#Go�7�#���޲2g��(t�?�!��q�C��%4c������]�S4D�j�s<��Q��gF�t'��g�Ӄŏɂ<�Є߂���b|�9�^{YL�B�R%4}���މ���$�ua�й��}��-U㵛^oD���X��A��ř�\m��(Y�H.{�셳��/��E�Wa"f�4E�l~��Dp̣�O]�	]3C�^u"ǹB'���y���I�7��M���3��+HO�MzD�brȞk 2�xm޹(���7�"�s٬6��I��g��$���tOҰ�����ԣ��D��.�uЧ���A.j�)��BƜ��<e.�p>L�����2;y��x������"K�$v�y��3-&�K��Y��&�60���%ϟ���0���Dm#�2૵�$�x�W�p�r俉�?qe��t�e�E��w?+j�˘�O<v�gR�x����J�X�v�&䌱�<�l��R�30X�T[��#\�~��4��	"�	C�/e�'���x�38WV�@]����5�f1Ǐ�`̎�o����k�5
�#w:9���@$R��B��B�n?%aw�V��9�	ø��7�!�O�g{�W��g	���\�ox�{F�Q����2..p�I4��o�d�"q y\4.�%��7���2���q4���<��
>�l)������k���%��d~���"�#B��2o�#9f=_{ɳ�#�L���/!�DU��OP��I�0S_��
��|��/v��ɟ~%K.����9�JԐ���Uq]a�򄾆�mw&��,G/���#��p�����0<P6 uQaBD��J�l��%�䏾@��7�E1���u=�Q�SH �|s����z���2S�i�h�_�I�=���*�_{�8c7���=c�s�X|�]j�cPA�Y�;���/���7?�h�g(>�$�'�64�pս���OO�.]��7Q>Q�Q���Q����+�b��4A0_J����KcI�`���c�}���K�/-w��6NW����O�x���\2��D�̷Q:b0
N;�w�>4��n�웈���eb�����'eGk�2'9k=
���4r��1$넭���_���9g���'t�������橿����m=˪�������`$��zP2
O�/)0tu�ot�r�Ng7�����t���p��}fuE�BU|4t&�Qk�̢����1��kK%�����`���\��A��sG���є�3YfҸ������1��UZ�z�����M�G���j��Z�z���%�����qw}xP߯�g+P��g&}r4��:�-�ݕ��`����6��),;�DV	�{�ϣ������H�G�[Q�'U�J�'�7S���[: qB���u�u4�WUw��0Ɛ�S(�2G��"!���0�o'$��3��?۳�&��쉲~=�#MLV^h����@&`!!�L�?�uI�_�������k(����Y�QG�-A�=c�g�?{ڝr �PY��迾.*ܧ�[WUW�Z�e�E��գ�Q�C�%��H���QE�Ͷ��t�(Bbu"F!`�M2���eZI���T���)�&*�Q0b��A�37�f	$�],;@Lt��S�̤�E�E�5��`�c��=B�7����XE�Շ�eE
y5]��u�H$,������|a�25�Ҹx3�*9�� u\&˜9��Γ�c۽Wmٞ�q���.m.�Bx� <b܄C"�Z�^��CG[z�`�^G��9)�s�0�l�`icY�8֔�_@Q�P�'�Cğ�pƄ)ڍO������joB�7�X٫��� ���H��8@�f�V�LZ�PC�����k���{� �9ƥR�Q�`�ON���?;�^��;^o6�����s�����x�q:�'�����ԛgص$�g����OA�e�����-���J��TJd����YL=�]���߷�`� �&K�
��r1O_,������xu�������gM�������.�����x���U����+VC��e\�7zȲ�C����	�*:�JPvNx�{��u�<��>�����yO�Q/�r+q�0-��>�%P��� ,*ˑ���b@���O����eǐ�y��O�tTIFmTX�9@���D�,�g����ܱ�Q=%d�������Qd�N��=ꍿ��싥ϣ��هoI�>� �#GC�㋊���e���x>r��w�&d��NJ=	�A���H�,���Q�u|w�! #�.¾Ȼ�|-��t	���UZ�୻�B��Q��K�n܉ʞ���z%�F���:��iM�3�]�=�9А��ֺ�l���Z.Kȭ��y�ndt��V]�`F�7^���?"�� ��>������ �R�^�+�|���ǲח=�ɏ!v�o�#�F&i7��:4���ͩ��O�:�ޙ-��������)%Cz�E7�XgK��_6�og�zB���H�e���	�qU�u�+�y2~�OQ)���^vޜ)��#�F�E�7?#ﬓ@:���y���\���z�ݲ��ֵW=z�\dp�M�mn9��j��ȷ`��n�C6~��<��%�}9��@�%�����;$���������#dE���������7?��>	kYz�1S�[�x>���AM�H1�U���ȃ��
��O�@��OE�%W���B�]�
��詎���r������I�����GF��!�~��+��.C5�6Fv�6�>4V&F���Qgw�񃂳��K�z���W��q�i�HL*y�b���|�{��(��E��w	1�8��;S�g/@�[�u#��'F��p��f�8	�zya���M4{���|Rc��7�d�>C� u�v�J��N�x��.��c9�I?�D\{�l���m���!��qH��9z}��%�R��ѧ+)�1���!�~�6�f��vb4 �k��A�E(&Q�t�.P�������%U�O���{፮!낷��������9m��_���%]o�O?��A}<D�q%e�#�e��+�����?�Fh%�Qw���y����^��2^}V��BV�q���O�(m���J��5^�����I���2�$�-k6����}+���+���@�p    IEND�B`�PK   6��Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   6��X�1.:�  )  /   images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.png�yeO�-�Bq����.Z(�����-,V(��Rdqw�Xq�w�E�J��H����yor��͝��I�L2�|��d��5U�	100��0%����?t���	��h�#7��'S��s�A_�?��K��K���������ח��孧���-���}�4��-p%}��c�4s�����ݹ��'N�"Ł�`my�׊��Da_����sY��]��`�~!�6F��	q�8�1"&��^��.=U��>������6�^�>1Z���� �Uw���I��1�vd�6ǐm�O�w�#T�7�<Bħ�O�Y�5��/l�8��)��*�ǥ����K���f�G�Dn,*��:��֘�ݜ���oN�`���쪰� �<)UjJ+��-ݞ=�T嬞o����B����0��p�W�	RC��r��",�¦��e��7���P�A�H�1��y�P,�F(�1}O���6ez�>�uby~���I��ڷ3��j��$<�洀H��%��;ϖ�o�V���$�=�+6��� �0����@s�	h'/?4�M�ίC݌ҕSp�u�~���-���x��귾3kF�&�>9�ڭa#|gTLw�ܟl�5�aI_z�߆f�~[%tQ5 ��:5���FjH��������fQU���Sז���_�8�w�:+ ��/ʦ+n�q��n��<�"��Ԑ~|���:�4�1=�ݡ�/'��^�E��8�t�f�x;;|*��ǌL����������4��?Ż)*�9�/��W���/.}�i�d͜���Ss72�6`I��3�������h������پ��I0�R��)#dg2�w �BP�p�N��	�
2�6�R�h���[��[�@�X��(��
O� ��A�޸�������A�m�	�Pn�*E�'��CC*c۱~1Қ"Y���k
�臨�RyL"W�x�E^��x\o�<>�|�z3 Is��$�[�I����*e�m�ȓX �рH)4oD��d
�X��/"d����h��q��}_W. �4H�$�H��E��k!+�k��~��x*{���Ģ��-���( ��h��(�|��7X]D��L��oۜ"I;ZCo
w���;��-kv�5���ID�Z�'䃨#z��[_IY .����S<_����cO[��u��^D����T�yc'�n��N��Y�C�h�ؓ��T��Ҳ���6-~�|j�������\����4�L��%-Q��ٔ�VZz�6��U�N��%Ď"j��\��!����u��I�l_�Q���w|{V��Ⱥ>��Š�����n3|x|��w��r2,p����m�W��s�I)�C��;���T���p��P�g8=�G�렶d��(��|�T����-��iķ�\�d�/w?Q����6��#O�?���ˈZ����c�\֍P�}0��G��۶Yhol���TC��F�%r'��l֮��o�x_���_����GP{0/�Z��Ӭ|F�L@a�.��s���|�3;�٦9���u�%z2=�9���wD�Z~"u�Nk��1y���5wϠE K�<�zzzB*������+��SR~����	G� �yw<QiG莆�������ʭ4�K�{��u���j��Ѩ�ft����q��42>V��CVo�!n�B�����=��!���_ʕ�c��'6��~��f%�k���&@��R��a�5�e��XDo�{n�̀}�wǐ0d����̓ �P�:������jӊͮ�!�Uu�7�Ќ�^o�S����܀��eI�s��|7%r�TK�������K�du1\a;ֳO!�Fz`E�����ބ-�����Uv�����TƳ.��]ܮؖ��.v�bA��.jM�Ǯ���������.��<���2��{r��""��Y���&1Z����׍���u#��G������o��UE�;�~ʰT^���]2*-�J������h8~�����s��:��~�l�h7�Wg�%�`�	_��U��:A��!3:iZ�^T�)��ʴ8Kw4\-�/��~;��e+��1Z�9\�ap�pb��leaE�]7�@s}t����X���� �Cf献/�[��u��kF��[���i�e�`��aS	mH���F�;ўH,�Q}C>�{��gذ|,��Ŗ�`
9�Ӫ
:P6���%� �84�H4G�b�},V���h�Bg�\[��"���0� �o�פ;*��Qv������p��3w�����J�#�G'Xq�i����"����Y��7]���T��'+8�9�$_V�TN��&�|�g���5�a$3����ܷx�fo`��܉?O�j���n����S��+�^rA�n1�b^��U�"(X�$���5��q1SH�J���Ʉ��$K�Qq/���NG�O0�h:�}y�[�.&j� �+�ma��yr���5��З�(����WF�&x&�4��[@9�ɪ�tmF�	����9�E��~�L��$*���\d�o����齬��߶��9�V��@�V�����'yG'X�R��M;�ˆ���%>/�$�� cv���T>��~�I_��~Z�Pv�޳_g�d�
U�/e�p͇����3�s�c�*Mi�!R�ث�8Y�	�N��YSud���d��y[�l����/XJ�v�)��������ٔϾ�fs��a��$�g��5R�����?V��-p�b����3��z'*�~wWe��F���9����W�B�_ZL A�,R�B��,zֲ]y��^ԺR���Y�z���D�J0I�"CA�����0u�]lC��j�� �Kr^!�������Tڸ�8���ϰ $,S����W�k�ì$*�3��,�0檋�K������j��/��s{�É� �	*̓�[|����nM;����3�+��V��G����<�0��4Z0�:G��Ps�Na�:�`U�z��������,đr@(6cV����N�ئP��l��;SE�6}��F���}[UC���v��Y�?6�j��\8�jabU�3�AD�?/��s#���7N���B�Cr�C)=^� 3.�_����1�c�1�t�I�9�t.�`4��
���M&q5�ޞ^J�Z+��1t��8ii(os#�6�(�g�=ϲ^:��Zc�����O��q
S�����!C�*�]]&mQ���%?"_* C�E��#�
��J!�F�]#�L�-s� A��c�t1s�[vn��qۢ6�.�cڶ���7��~jJ��:z�6�A�?B)�լ��c���n�U��ceII-�t���Y#*������Kuv�:�x�<�S�h/\�C@�Ο��˝��9Z_ز"�o�� �Z��].�9�ɵ�/�W����"jQ-�0�+UOQw��8%�ERV�.EbM�J���b��[�AA�&�Xw���5�C����B{�"����R7���$c�R�13���?.�T hS��e٬H�e���̱�*��Ҥ0�D7��(TC_�K��&b�	����zX����>}C��}$c-Ag�H=gwٰz����4V��MRp��ޞ��B�������lyyb6d�`��I��E�d�K�q]p�d��$��U�H�L���D��� �MY���Z�����*��CN���J�[��5KK&�����Q.4���������Kk��U�t,m^}hg�p���^ϻ���Y�6-�ݓ2:N�i��{QK1�@C=�0z�Az�=�PL!´��G.~�:	@��*�{��r�d��%^)�����������/���Ո|�b�_�n�d�'%�%�|��_m��zKW�#�Cͨ��9����I8d�봍��rS9�ʚ<gX��a��z��+�Q��|�l�,+�����U���ƉP�B�Ix����uX��с桨�y�q)>M6[�d� _q02}����IV1��Z�YzVw�|*������\E9L�%|��&���OI^/���P��'�q�M)y���(o�F�����A�3�^(~n��3��¢�Mbt�Q�0��[{�	��@�8���Յ�^�e��5�>j���^�@iI����w�w͜jG�RB���,���qK�qK��_q3�c�	!=uoGi�,���EA4�kk��=ҢB�}R�e�\�ቀ�]��[b�������)�j���#�&�4.�uu-�!�-�T�2��i&ig��p����������	ҙ?VA�Y��^NcU(x��J��ѱ͏p��ص�sf:��3^~#�=2ܲI?���嬸d��xN,��ΤL@���rl��z� *�Pmq#����__7 ��H�B<j'r���I��m�H�3��\�hxi�[�q�ӗ@[,������%����b]�pvR��Q{��̜�޵뤗_2�)y��ѝ,km�R;D����2]�L��R������n�h�9|X�q��a|i�
�W"|6^p�[�Wȳ�븅�`<kN�Ә���?G5�^l��2O�V��]7	��0��m�:���PY���&�%	'j"��,3cj_Ns���+`qA0


M�z�ax�(�)Ƀ<g�5$�0,�t�<�1ֽ���lj(�`/#�g��}���	,�}���8F�&�b
UQ��!;�b�#b'���dV����@f�(���\���S����#h��O�:ݼ��a�XVR}i�һ\`��\`��D�m�K=���}�ITw5!��	���
~�n`()xz=s�3�.B�f�X�i�k�%P=�Ԋ)�jcɶ@��q>t�M}�K�/xW��Iuk�[90��o�A��dy0*�I
0�Ά���}3�?�O�V�m����|4(�e�OӖ.��-Ɨ�����<��ϱ�#E��x���i`C+�D��+൐��T�������1r �^NI�i&c�u	_����xi~��j�o�t�>�d�S��,%��Xd�z�7i���C�_�{���⢫tA@z�.�S�}4%Ь*,�{�4����Dȩ��L�I���%K��g�%q���w�y�_�c�{qʺ�L0n"/�����zt�/0nGt��d��G�=�x�%;9����=�б����&�}�+�m��s_�l�bV��S��;�r�9�.W�i�����F-;6uoN��I�l��i��~C�"�p8�C�� ��؎�הݮ���%���l���ܕ��1k�:�g����=���{������G͈ne���$�(���^�������q���[�N
���D�h*��(�#Oht�aq�|*�t4E9��mK��(T���]a����8���f'��)��z��������\�t)���'�����`05�t>���Mt�=8mx�U��&��@F�<�)�^|�8� ��w5�j'�=�M�w[�� ���&�⸥��n��Ǧn�!��~a����y�
/����'��ڑ�9dW�����2¾5��.�#�쪩͋�@Um���ZlK`v,�]�#�>�7�1�a�d'�#��F\1�c󱢙�5��i]) ^�8PHN�=�"�D1��ǥ����аf��_3I
�G�$"8�0%����������������[�!���8r�kB/��S5c@B�ND��|�X�2��v,����\�)a�]���d:0N�s����o��\��ʈ��Ҥ�!Iu؆Vs��*X�tq�֗}Ȩ\��a��n�ћ>�Vt�ye����w4�F�)����n��oW��y���V��D�e�(/N�#]`z'�`P��ec�����H�Ħt�����O�]��B:�S����I�a@)5�J�z�@�%��9���Y���\�+���)��M���
J
G��y\�Z1'�Xߌ;���T����yS8����:j�!0-a�H<8���f�$��i+ç�t���!>�A-��\���ϵ�� ;��3��4o�u�Iw9f���f�4"�h�m�$H!{�O�g�c��C�C�)��ঢ�S��"5<���3�o�9���fK�!.�������f�^M�Y���T&۴Js����n�"��B�|�o�[�9l`���2ˏ��WC5���-�Z�C���c�zo���=^t$�[&ˑ䨤}�JzgM집D珦=o�M�[N��p��2�u�kx���ڌ�Ȱ��y�+��.�T2-�SJt�-�k��]��.��0zX�h
��ڒs�%�E��>�e��;��ã�/fMۅ�]j$8� LA����F�TM	��{|��EWՅӀ��"�õ���y$6 N��jC�^�&^k�DL�Л鴯SD�i�yr�,?PC�b�^����N�y�P�tm���� w�~�/q㵏���&����Uq�б%@������� �U;��?oT�-�S��4�j����JX�/���yH��v��Iĥڰd}f�kه[�[eo~i6�y+[�2�Pw�2Md��7"a	L�I!$����GNqZ�m�8qI{���;Y��l]�u���������Yʖ+��_��y
�.�h��f7z�\U���}�S"�y,�fP�Q9���5XeYL��?�.�������]���+�Z��9�j���,�S��~���:�=��������t��P����E����@tuX{V8z?Ѕr���k����7����+9�����뢓oC��f,�QM����E�-��M}��r��$����:�v˝�G�4�]Bp)���q��-�o>�����*֏���ץ�R��-�rc\'���F<�"������\t �$m��@p$���]-8�	Ǜ�&����u56CӐ�Q�� o��j�}||}Lk�ů�H˓��W緽 �.z���l�p��drB�1-E�� �G���v#q�߆�[��׿_A����h@f {,��ӤB�0�B�+9@���ȉ����2%]<�Ǜ�9����ɤ�޻��
"+�s5��I���N�t�{+HI�~���Vr��� �D��v<;�n��S<�x�4�at(�B!�n�#��J;�������>�Z˔z���L���:s�	����8���8<4 /���q���>�5���^�P�1�C0˓��2o�y�����o�Q�,VfϞ�իwCR�{�ϐʃo��*�� N�Z�+'M.��mݏr�)����(u`�{�e�M��9|����/GD=/���BJ9��.���{�f���������(��5a�vx�&�V��<䒛4���I��6�K��e�/j�k�Z�s�2+u^�����Xf˻��{k���s��ZY|u�F z}R#��O�:�S_�E�����ho�lW�;�T:��z�K��і.� ����mjr�b��lT:�˒�:T����Q?�y_��_C���]�3�^�I��.�$t��@��K|>��+�%�;&`�1�έ��9�s�@�TN�_&C~ͪp�Z����
HwTS��L�Pq�0;m�i�4�w{,X��+�� ��$�uԡ��ۧ�~{�Y>	#E;�D�YUq�.%�[��E��S�V���R��n
��O��:t�m�D�6TѪh���lF�J�ُڇ��Ev󧟿�
���/�������\N��#�_ J�Za���/�J�κ��Ȕ��w�QI��dˢ������j�%a�dP&���GW��W5v����n$h'Z�r��Q����R�.W?�MW� �Y󜖱���A��S�_��%=x *;��f�eA��y��#&�}�>`�k<+�z&�x���AC2٩���}ŽQ}ָ`��{�T���+�:�Q���}+e��T?P���L�"t��	����-T���hf�[KzGd��Rʦ��7�Ü?��	dX`M�-V]z�#��k�����5�>C-C�PK   6��X�Ƚ׌  �  /   images/9185dcb2-65ea-4de0-8d42-42cedb1b5634.png�x��PNG

   IHDR   d   -   X���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��\�o��ݙ�����uڗ��!Q�Bp�D"��h(U�$B�F_���?�C�JM�!-�А�J�(�U(I��E�|�^$k�w��u{�ݝ���?���gM|}?~3���眹3'֎_�A`$�M!p�8	Q����~��Ql18���gv`��ű�K�Vr���x�p�z�3���rW�y�4�0Ɲ��t��=�r�Ҙ�xq�!4q]&��:׸:/s����Թn�?V̕%�p���:�+3xg�X�@?��Ⱥ�qO�W�t�G�����X�ѳo���Ij��;m�I�Ae�ŰĠaä���	.���'�eV�	C	��h�*��2�z�=.�q�k��I�%WZ�A�KD����rB����'H)��8�{?J����>�9���v�4�'���~��.��7�'`��9F+ o	�'�!p��/e��!i{?�CP����Ij�Ҹ<즺aj;C}��Ǘsݥ��N\₱�ߧ�$ސK�\��G��	y��s���׸��s��%\�I��,� ^�cg���CT���;s���/��e����2f�f�}x;����Q���r�����2	��b�\͘�#���-��pb�w��u6�S��;92���&�}�5L|�,�a��ʚ�K��D1p�eM�H��ugDq�ߣ�[5.W�z�D
!����	q��MB\s%��Zs9ߦ{�/�$��b	ӓ9����M%wk|ao��3�=�)㭱�I��4Me����K�_�%?�q�<��5'��-����Ү_���W��:�of?�˸S@�w�ۻ��~Ϋ�1\��K�
�^=e4��"������W]�r�\�ո�k��書��հÛ�����$����ǰS6�}�������>��ذ�)���Ty�"��])����ZMtXT^��s�V>�q�<C%C�u�2�~󘫕���M5�;s���R^����D����}�s_!�.I��VH����k!�){a���2��0ڔ[���̵��`@��XxL�zp�f�S�7B��"s���q�<σ���ҿ�P��J��h��Ȝ���g.����U�^}Qx��t:��C�Z%�d)�jдЛ�s�1�J!�H F����R�����Ӓ뺈q��U!�M�#���c��"(�Bt��]R*��V }�����H'��t��Q!���xUH~&a�����!١;غ5 CG�4�O4䏱z��אi4)D�Ζ)�L�8:$�U�vQ������:�Gx��x�.��~���n#���q�EA/W�W�H��s��������/�]]T<���}t��.��j�G�E��WX�_�|BE�
���Y�0��/-S���F�]̓����@�1����n���~k��j�ل�C�ޠهđ��CW�c�+��+���\�B��T����8���u<6:.��aYC[q��Z]C�r��X	�z�Z�Z!�Fcr=�/��Ut���q�@�\Ѱ���\�d�\���r�r>jp������!�=w��B��B����`t{c��	��겻�GA��lZ��v}�m��_�Z��v�qb����/�^�B(JKO���'a��iw4���������~zHي+ڮ���E�S>��W󉞻�S*;e�d��vr�-�+�hVXG���f䫊u�S�#�J��Uj�pc��mw|}���l� i�!�x_~=����oܺ*�5��S������q�8N��\����MW;t}c844��'G5���!����}yB����a9F{(?"�_�$9�c�3TC!���
)|�B�O����ؗ��0�W&�RxT�R����s%v�iѥ)��	^�U��=+���0-zJ(���/����R	o|�6��}� �3n�����=zw�G�X�ξ���z0;���<w����4^y� Ο��R�¬����i�C�8��y,U�0��UI�c��W�1��u�Q��\�����p�{`�OO�0Br��V�u�0���\�=�r�9=�Va2^��ͅ	!�sZ4+���w�n������ة�jep��!b�~?�7�՟�{PiѤ ��?�(�*��    IEND�B`�PK   6��X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   6��X?S��� 2� /   images/99226213-8268-43da-ade8-d9d07cfcec9f.png�gP�Y�6�3�3
(���J�80�d$g��AR��!I�,y�$9i����LJ݄&������y���s��rW98���k�u�k]k�C���.�\B d2O�VA H���$��̓�_~u��Q#�7��+��w|��@�� ���f��
|󆋔�������DrX��8�<w4�pp�Hŉ� �2��架������ge8p����9~�����9~�����9~�����9����D�a �6a����s�?���s�?���s�?���s��W��
?���|���t�+�p�����q��ds���,�r3�A���7��vaj�(��%'�	�ψk���XRKj�^ی�����~��Gz�޼nq�"�s�lz�c��*'��B���G��*����'�t�����Ð����9~�����9~���Fy\G!�~���AN{�8�֤�M�,�-�U���0/��w�Dd�-�h/j�`��z���L��qe%eP�Td6�`�$!{+m��+�H�0/0�EV\&.1����2wV�6Rer��t��=	���n8X|��^�V����ϕ���-¯%> 6#�
{q�$-��6ﺴGDW`�3�O�5wr�~�;�VNYv���.�7N''kg���}��:�w4&vy
|�4;�k��:�[�$���L�Su��u�w�4���Yz�+�,$d1<�nە��f�=*�����o-;+�s߾k9�����#����0I3��\�#n�-�1�i2E�=�]KeS�g�~Q���z?K\���N}��N.'�M��x)~M�銶w�����2�-#�z!C�܁�����k�U�<K���5,Oz-�e"l�k�xͦ�ٻ��Ǐ�U2�+u�D��uLǭ?U����{3Go}�5$H��67�Ck�g0܆�����<�s���?H�&�����i��rJ=��k���p��ҁ�Ɇ߿Q!aYP+ڭ�ұc�����X�."ί�b��$��f�@�ى�a>�[O��w ��[� _7+�����~g�EG�+�}X��$�qf��q�VB�<��C�����B�o����Y�xj������g�bh����>�ޓ�̧NLPK���ߨq�nd�����B�[F,���O����o��)<�j3����J�-�}^3�S����q�o�'<}'�0M�F��`7�bqmwi���~3��քQ���dFK[XQ�����5����b&��-wd����^H8c�V�g=m$�,�l~��"\D������ӕ-��/Cny6�*�)�O�|�����8�??~ZK��ɳ����[rm�2�#i_j>���1wY��l�[8W.5���P��D#熆�L<������"����Q]��]s��蕄\�y"���;�˰��G�v$��T��Zۭ*H_ݥ��<�>�e�g���P~8FoY"4���i�ɚ
�29�
��g�'٘,�����%|�}��ݙ�F�k&�{ټ
/���\�.���� B�v�ώwt�m.���v���2Ln�E;�3&�e��Y�zDU0�GѷX��R�޺f�&�]0x�;S��>	,	M;R�v�-�)�Z?3����Q��Hs��H����
�y�٩3摝je��4���%{c��E�[::4j���T�/��~)0���o lC�{�݌$O�4{!0uUe���1c6�s��a]�Z�~{0�X�����,��M�4-�F���z����;�N<"O�?�4�q��|�ɗ��Z�+у���[��*�������^�Q7�~����w�㔭�S'����:�X�,�����������K�b/~0
آ����nXn��z><Sj*<�Ij���}{��J��⃖��.���C�\�r�J�l��2�|�-5��u�I�>6k:��y`޸?-3��׺8;K�{�H��d���A���G˝�����ȩ>�ZhO4�h!5n]b�ݫ���R�4�W<+�Ej��7i��BS9n��;xZ%�	?�8 s�<n�%̝oz���(��-��J��/��jX7Z�����(i �_N��Z�û����y�soձ1w�7������2UOZH�N�-�Z�G�(6���oEuE'�pu0�*�S?�=_B����"�/FW=����ټ�*x'D}�}�6�
�����u�:�j��:�lГH7���3Hk��?V{�X�pEn9p�-g1���a �������5��!S'�[ԗ��<`uy��mZ����ݣ�<n�LKǳb��c��`Y�4=�t��?�����>n�~=�-?�1	�/s`|��R���x�g��i[k�����h����__�J�U:ڀ�z�L܃��._{�(�%'^�� �N�c�e�ڔ>���©��3p�B;�,����L�:6h�z���"�Qy�*��hu7r+�Z���y�6��s���Rv����Մ��eܹn���Y�ۏ&�>��[M�L�T	8��J��q>�x�%�ɦ�lx;��ƙY� �ZR�pf�u=wR>�:	��l\�����������(����`!�x����s�Z5� _*�ȩ��@�a�=v�0]��0�-�7�;��ձ�i�&�6_���<�Ik+����>fͨ��ѵ�N0CBK��R��J���j�u�X�N����{���R�6��t����`�g	nK�3rT]ݝ��B��6�|1��`Ba����9Ob9o4Bz�5b�V>3�s� �8	�c{7?�� ύ�b��.�l�*_����N�6�~?y���nTy�/~�8,'i<#��Q�n)��������h��ܖ���7��}��c�:z{��$6N�����:���g7ŎU4���4�}	M�M��f�5�����S��+��pz�e�� 9��BEؑ��#�*@hL�N��o���M'���E�e��h��$����0!���d����}) n�+�~�D�is�=`x�� ���q��$ bƱb��4���/9�0��������`6�������e-w��俀��� Ä1Koc�r�o�v�T"5>������?v� @(zP,{��9�/Yw9f�k�:ͭ�V��H�}��9�Y�o9Z�t��=� ��q ���[}�0
)���|���� X�E�������ѵ������M���Av, +J�X�<>��zFk`jF!(o�ӻ�U_;�����6}�`�p�=�5��e��������؊w���ǡ�����&����'W�Yɚ�HI�:r�������������Իk�oR�k�[	lJXN(a݃���-�������_<V��(��Ow�f�b��g~���ٗ�޷o�h��j�����铆�R�+k���)E��0�GwU׫��<�ݹ���Yh���.Gu>gx��l/���u��j�$y��h�����S�gE D������i@�V,�(��8,=be)���]i_Q�˸��|�FO�������1��U\�>ơ6t,��<;]�i���C�&?z~>%f����V�_���x�f+�,�`�����A`%���Iك~�llZ(/4��\g*�}�~�a]#�1�IK�
�o�z��bAz����P���}ε��1IŠEUUt��1:���0�{Ӿb�=�N��@��[������^4�7r�?H8qpߺ�yZ������s����~�y.�~�y�h� ���!~�2���0�����a&P�so�!l�;qp5	�RPW�hN�>���Bad4ڴ�h4�%ho��r�Ǔ~�}��ܼA������~NGǉi�_x��	C�����  �n"���P��;�Y�th�ԉ����M�!s��y[�y� ��2ǬK���CKF�4�f���ɾ
/��Ryp�`���t���!3��z�{F�Q\�[o�h�(�A��&@�h�*��E����U\��Hvѫ��Qx��0W���z��7!��$t��2���,�mO�����xj�ǋ���p��q=��_��7j�
���S� b��o����@�[�_j��(o8Z�W1 ?"�4#��ɉ	�)�Y��E��<��f>͝�M(-���}����E]u����&�j>��b�}�h�`�r��*� ���~�
dG[���s����'{k�����hvPO��L��_����/z��O�	��wK�D0�P\R����=S*���Mx�vh1C�cܑ��U������z �
 ���Wx����ܽ��aGn�s
��P� �����@���Z1��{x���+.~0>�[ ���큖Ԝ�jWGwynˏYC���ì+��֎������<����jEmX^�J�����d!�kEE-��������A~QD8F���İw�&~�p.��B�� jͬx��� q��E2�@S���Z� q�1sv�t���+,m�@���l~�5{�R|��� U@|��40?��m������F�O��f���:���pi��+0G����$`�ׂ��g���Ϋ���>R�Y�U_���om�MT�xy���]��;=;+�� %Y0fqiCܱ�>A����V�<��P��3�7�mf��w����pg��j�@�i���a��R|�R�0����hh�2�����_w��f����������Oq
A�j�a{l��������}PB�~`w�>��&��(��R}þ�E����o�9�X m%�s+�F�����ڽ���%q`�y���S����9�$����i/F0U��g{���O=�٣�;�^a��SBR�pt�cݛ �d���[����ef9�KA�v
��\��|�̜$�JN��N~u|�k���\�6�d�/�1fTpxog�2���?���'0]��z_[hId�߯:K!\����%8����}|/��FV ��((�~��rV�ӓʏ�x1�A�ܪq�ַ��Ԕy����� J��R�eT��m�~�ǡl����D8��\ЃY���}����;9��}�rR�ܷRR	3ƒmͧ{��8� �(��*��XD��b��2K��z�
���ݵuK˃�)�Qî~ȩ�PNh���M�,)e4��+����gp�X.xtd"��U�gS�xmخ���%Ey����ۇ����ع�����)c@��r�?{�TlH���Fn�U8CFf���������!w��|#���(p�7�x�b��6�ii��}6����b��?tG��g�K�R3+�or� ?d�G^��2�e'}5��Yb���s��+�_������5��ܤDV9�P�ׯ����^�

��3��ׄ!Tφ@A{5�E]S_EP��GH�l��%��a�y� ��#���L��RT�-�X2$ز�L�ҧg��Z9m���D�\�J�+�rO�ijJ����I>-��y֕R��1�#��s��j�"�饻�FoP��9�*e�F��{}O&vd�ؖ���] ���<a�%'���FFJ|#(��\���-���XcU
�{m�.|�Fn��@���:`;��߂!�:�$��I��-����{�	�+BQ*%O{��N��d}��K	�����(��r�������}��`���6B'��rV�FYv�w-u��adх����ވ}F:&9"R?��@];�X���rb�SW��>��'h���Us��M6��i!Q��oS{9ʖ������?,rUPȴ_YK��Q�QZ�����ҽ��d�cc	2��]�ZZ*		�q��^�k#>�xlE'�
��TyN�����_�?[U�ЄL|�ܷ�����Рd��1C�^�J ��8�(#77��W��1�G�`"H�^os�>������_M}WW!�ӗ�֫���Q��1�Y�gUl9�_=$Z�,�XJ���Bh�>P7hM�$)~JF&=��(���`=���ֈN2��8:8`���_�v�xˁ���]RD�;;;�����bL8ʇ���^�N��[X�����d\�DaC#�:Ϝ����Z_��{t�w���I`u.@f�9J���Q�jk�?G[�܃�»�49]�����­��Nc��FCO�]��I A0�N;i<����KV6k�$��%�.�<���:��==������*��pGx\-�w��G��v�fE�#%2TTb�����7������A1M������ڊ�ܗPE���͈]?�'��B��hg_{ܓ67��V6��/߃\^��� >��zm�D9�̮]Y�3K������?f�f��9Ɠ��-��M~g���_5�l-#� 4���lA��ʸհdc�m2��h��"��ۛ�)�j������z)<�>'��)��K�anD	U�_A�g5�!8W �F	g���'MZM�vy��@���5"���9I�/0�;ux۬�.����A�N�*Ha��46�M��<90�QZ���_��k����y��mv
MoO��t��ׯ�+�˼?R���w7&&���\��}W��2�
�E
�I�Y���zC�Vq8�VO��z:III�+/��v���|y�}�.�2(u�٭[�~:L<�R��%��5����$�&�f d�@}����A�q���~��a"��b߬f�+K�U��S��t"��LU���Ch����2Y����:xP7�op��ܑ����?��k���$~6RH|(v3��7�~��s����0u��8D�T�M�Q=��7����}����ct��is����F�\��h�_xG�u�<07W&+�H 6�ZI9T�V[-��8��kO���"@��(�LN=���C3zCqPgHb�+)1�\�輏����}�>��v��0~ܚK
rzg��%%>�f7*2==�i�N�8\��5���?;M0���Wa�B�_u_M�/Xgm{�^]���<�<���ֻy��綩.�g-��R����oH����? � 4����j�I�l�����8���1����m�\T�q>�gk�01-1[����������z��%(����s^�d}�<=�����8`��XPK)��O�GEP�,�A���/��mis��;���k#=��E/�]lJMO�̮�0��m(�uA��:%���;��I��o=��0Fo����7��������� @�t��Vx�,��g&����<��.d���yVOSRn�Jk))�'�cHS�{�r����u��&[�{=���3WI��.�`D񵋬 p��'']��WM���kyz!n-|��E���^�sJ�X��.%���NP6�h-c�(���$mm�qY���ujj�е�������1f.i �[ix������N���1	�����v�w�c\GO���0̟w�)rߙ���W8�M�������:)�q��- �s ÈL��V�?J[��Ɛ-��蘘��'u�ZxV�1���c�Ų��t���3�e9�J��� ���*k�,���pt���:�
h#,|�v�r�[[3$qq�]��}��\�n����oԋ�pT�A�対��]�f�5A,&"�a`>S�!������x�!��w�uX�&�@vq��5sߠ=v|��� "l��q|_�[�?^�Tt�1fخ��K���Jyh�@$����<
��,|ji}�������F�`�^⯰��w������H�A1tt�+}c?V��Q?��'px7X�5ޕ�h�o��DN2~�8��2%%4��������f�A����i�!(��
u $��SR��tt|�����C�!�Z@/�o+�{�i���hbR&'�(
�e��қ�1�̋\S��$9#J���*�:��P�J�P��\�h��\�2�u�Jaa^lT�.�p�a�� )���f4����W��ǝ�� L���ό�z� ˤM`rI�?o�XWg��}����Ȕ���"��'�3��VT�kZzh�Ǟ�.ZP,�_��U�ЧOd2Y_�C���jh�f���z��!䏆�}�nI������P�#Z{(c���������b0�@�bv{go�8?��~DD�ݾ�Bx�,ϴS]\�_�M7�w)Bk�MV������=>	�����ק���6)�q����o�����v{�Lg'����Xk�
�����?�ne8��M�K�n��Dw&9"�LBK�2Bc1;�ާ���ʐ��3t0ם�B��n@e�**`�RS<�A<o��$�����1����W�I;��V�_�pp�((�ο{�A�w�6B&���ق���V�����*�Бf�]w���♹�0���V��f��jN��:�z��Ʉ�Z��m��l<���_���X�^���ʰ�o�Txl�Vj�-`���xg��ηe��8�����m]�@���6�_����Ԕ>lb���mH�hV[�44���Ԅ�)R�y���L7�܂��(�w�A��bP�T��b[*^dL��+烲��ꊠ���̟\���C�&&W��RdL��Í��0�F��uV]{9 �^V�~~-��E:�
Sz\]N�G3D}�,�jkڬ���Z�?qssu����0{j�(e.N�����a�`�+?���:�R��cN�����g���,~���FQ8�io%G����u9��F8�h9����е��Y�t��qպ
5��c5���S��oߐ�a��J'>�i��Q��jZ{�"&�j,����|�������@g�����K��%����$PZ��lE��Q��O��M�`�(�����11���}��4�V��0�x �s?jC~�E���*�@tԙާJX� Xu�:��=�:���΍��X&���s_nnL�R>�XB�,~�r��Iw-�����O$�6�h�ր��Q��F�皺�)�}�ߟ���������-Q?yr�P���X���51��Мm�u��#ynh�V�Ųk���c͆៌���4���x&��Dz0�G⳰��q��I]]�T��F%� (��N׷Dh�hB��<����h����\

�)OQ�s��������LK�ӣ��p/pL�&�U��V]�m�� ��a�� �S4M�[˓��4��8KT*�4g�U�=��s+&*�Ã-6Z����6mw��(����Oc��n��89y��'$AN��������7q���;��T� #��c����V�/ϟ3�3>h���Ş���#7�{+���_��� ,rjKv�wP8�_jjR��kI���K C���I��z��Z(��wuq�gap��G$-A�I��c���śx���@��׵u��Ζ�^%8)o�K�L��`�z"#O}��Go��)\�li�[�����Y
��Xik��JFn��--7�5����E��pt��]_w�Q�~NT�^)�w�'��؄K�� b��h��j]���͖0���=��Hv9���K6a��k�K����4�j��JKҪ,����eg����s�y�����Ѡ;�ɨ�'�z�i�x����0nϛ��b!�l���-m/�.���D��2CBs'X#�X��;���p�Ç����BIC�9kXY���˝z�M�JI�xQv��D����5�T�[IA�%:���B�l�A�F����A]!�zNR71���R�������z��*M�.O_��Ћ@��im5������h�jg�e
?6f�5�Ɓ�m��������}�$��#�r�Jˎk�]_~����WRD��g{��wvFs���㷁 �|��!mk��/���0Җ��q"��E��G�3�Jx8n�+��_�N�uaH�4��ڕi/�[0�T��&A�S� �0�GR2S�܂bKE�6�t�~=j�%P�90+Kek��tHH��"qyy�.n�K'��YpG�F�b"@ߊ߸y�#��{=�k,�']E�ȴPe���"�������h+�.���"q8�-�7n�fXXZ_��y"mHZ+�����L��vF�5g{�Q)�ʤK67?�%���%(9�i��?/�B������3���А
R��S��)#�����m�^\҅|9�X�{_�P[�ۉӒ��Z|�U5w=�1l|0;����/W�c>؞�-M����7*"n�M��h�T�1�,.r2r��/�X�Ud?*)��P��S��'  ����~��e4ZI�e�������h����sIL�5@1�y�p��6��l�;�K��ixu7���߉t�*,tbz,�D�d/]A�n��&Y��\��\��)G�e��Eʏ�2V��c[�U]�����ڭG-�,(ߺ�D}��,�"�2+�����BMM�x۱͗@oM�		�ٯ`�����-�IK;i25�_����;�(_��u�f�dѵB81u;������p�CY��9jN­wH��1 Z���|Z�O��@�L
��q��x(4����h�p���,"qgU���u ��9��h��~`g?�T[ۜ5�P��< ���/���d�*�u˿C���?��gW����^��q/����\9��HJG�;��ejlx�		0DF2X\�p��Z4�e��
��Ϯ�L�_bT4� �h�$��l9�X�*�B��И�
*�Е�į�8�fnvvН�Cz�-=lI$���dm����{�e��M�
�M#f�k��X��p�z�x/�u.8g�
�����AIO!)��T�č�Zff��y'��܁D'�x⋲���iQZ^u����������sq�	�Ѕ�v|�wr���M0r;�(��}�����z�:K|Hp%k�[� �;q�|�1�>.]\�$4t|תʲַBSh�vXL���b��Ћ���\ˊJ<��
M�ſ-����>��3	ڞϩne&�������i>ܛ$>CfP��d�_��Q���Z@�s�?�����Dc*F�[k�.\�{hx7���u��:�l�+����i0�qK���(���v�3�4W���N�I
�M����]]�=�M��"�`ՙ���b<^�86F���j�*��r�N�Ec^;�����(���Տ]����<�#Ǒ��;���n�&2j��V�5gKc��Á�(̇�[t���T7���2F`.d�/���ė�O�a�	1j��>�L�}s6�mss��F|����i���Q��1r�( >����g��鍉/�'.�;T������2`ND��)�(�eF~(4T��L/?YHIq��p�6Y'W��$�{]���ϯ��`�#G�Ǎx���2�m��!��~�9�r��҆�թ�MFɬ/P�i�����bԨ Uj**�����_u}��ыJ����>F�4{�)9}��P����4����ќ:�����X#�]1�CR�wa�UW�-z;3����|"i@_��DI���Xr��B��U�B��.����;�z�;��A~�ݷK��%i�6���T8�����:X��x�=��4�i��Q?�Bݬ|�>�@��h���֭3ۆ�/�i�ߦ�_�>hR�H��'>�W��XK˛k�ܮ��ZZ����������X�5��2�k�vq�$b�e�"Ū��l��PUG{c��l�k�Cӊ {� ��n�4J(*L�vu;�^�G���Zd�" 8.9x��V���FD�C-���j�C�@&��l��J�M*+5��k�9�i�.�e<�!QQe��;C�h}ԉX^/�E��ep��E)��G~�j�n��j6�����O}̎��San�q����O�$�
(o6#.zz�����bNX��[���M�l�ll�@���s|i|ӑ
E<kKZS�M��ׄ��<36�[�O \�Lf�X�h����_C�_���X&��,��ǒ�.�FƛOa���a�{�OU1/���7�@{x�OSAM�Q��w`�����5�k�AA�J������>!�4�qF7��$� ���t
Ž����)�_�� �܃+k�q�='��R4�kr���	^m��[5�,
�|��3/��#�E��wI8表~��1���.�(�'67���
�}v+#�J��S��Ђ��0��z����T��g	�\��?���{��x;��V@g*��1���`�dC��k3�J���CG�$a�'�Z]�����Eig��P�>JRP~������.��QM���|��fa@��Ȼ>^Y�6����� a�&'�����[���p[��"�Q�7+{�ui�kC�|6袵��Lm1��P�⶗e섆׸Y%��* !_D0���/�oZZ� ��]N���Jq�e�Ǹ�k����Zi��b|���:;-/�O����������]�^����DA��?�V�����d~~q���¢�t;R�-�`��%y����QH���.�qʌ���6�鋵.3EG%^��c���$������O%$,^�1�!
�T"x/ܟ��ΞYT����; '��hJ���#%�8�]@�G�j0��82�+%2��U����h�˴�@>L�lĠ��m�0��T���B�}�6�ݕ��@����ԙ�k���m!r2$��������k��0:L�B�����A&`t��sV���l7 .�_��*��"I�+M���N����&j~��ϫ+CT	V�����F	BN	�@8��S0N��)���<�h?	`��[ b@x�>,����_=���	v�1x��e&���k�}�_Y^�b p�*�g}l����y������,@zl�9p���D�'&�$�&	;�gxه����:��NWAD^��!��wMG�Ga���̇�x2��K��X�f�� "ˣ ii��[�-O�M,pB�e��F+ˋ���Ê
�����P$5��N�v�U:U�['�}ț@��e�����+\Ζ��wL><j��A����tt�A �<��<��6��a#}�۬�3(�-+�ҷ������kkׄ��)�O�lA��NMk&�͓\���L%H��k���=9��u��O]YQH��ڠ��d=�%b�a��r8��(�N2<u�\n��J�{���� ���`W�Mn![:<��^�IlW��w`�'��ޏf�wu�^�g�0�w���(�3:���p�iy07�	��Z5CO+��^C��("�7������DS�:	�Q�Z=n���$l����E0�(lʰ�44����P���-k|�v/ņ��Z��)��Cl���f	�!:-ϒ�}ך�����m��M.�׀vJ���V� �g��������O��I�t��cq��\�fIHI�q�����-I�c�#��4�4v@�_�+*��A'z���fK<�k�a�{.)�N.�0S��1iP������@��<��Z��u"�pӧXX'Z�e���,$�]q�L�Rݥ�V�u��[7[`I�\i}��#��$FF2��\���K�`����N��xp*.*��w7����?}"]�0��X8�+�{�t�<{�,F�t`��l]Mʳ��?��Dm������M�<�
֮h�<��>���_R$G;}<�َ�ш~M'���}���}yAi�,׊FBw�I�̣��e��O
��VL�m��Q�����'-~dS�N��t��uOο
��j���r!�	���t'�7�}N]�GU�����o�7��mnZ�W�����2���3���%���ʭ[��s����L@�h�)��͌��[�>�O^�1�!��AI`�9!��d _�[��V�s��_'ײp`,gc�礯/,�kğ7d�=�%���OC�K�����蕾�$���w��sUnѰ�{�S�)ނ}�x����8j��|�;���a,)�m�m����I)�=1X��N��������%�=�5�<�B'�b𣞫 �*����H�
6l���G����#��8�Y�x��h���9MQ�Q �D'�Q�~R��?�ctW�b^v }	k�9����Çɾ���{J���A'�G������|J�y'w������W�_贮��(h����`g	)(��.���
ߏ�Y[.�v�����	��~4���$%K��ߡ���y�,
�k�/�ΩU��ԍ���-�MA��gB�U ��*���
�Z[�$����*z�	���g��������@d!�s:�9J�Xٛ�����R#�S"@S���E_�n��+��NH\Gt3���z��ʧL��r��q�Qt� zj�u�=�:�&�6|��f�J�֑��(��{��PuM�w�ѯ2�(��8s�W�py��	�$	�ߴ>��Z�b��Ǹ��*@z<*�����rr����x�^7t��<��Q�}�/��)��o����]�q[�7Wl�����Z/{
���F��{��[_J��>  �#�N�%$����C�#��*JI5�/�w�K³���;	��mp~��#H�If�꿠���P���|��4�TUf�'@�T�mI�3|���(��Gu�������4Y��7�����&0H'�n����H�]Mqz��,
���Q�IuQ��@,�C,V�e��W���JȾTT=�b��@� �FQ�};�����Zd������Kqv��-L��$}�w���2V��_���4/{�aRC��xYZ��X�%�q����J�ͳ�!1GM���K�*F��I��;Y���2�i)N"����둯9`�g�݃/-f{�T�}�����hj��U)Wע�JK�lN��ᗾ5m��A�)x+�#[ڏ�����#���5٠'�����_�9Վ3>x����O`()5X^��t�g~E=��s��l��p[�"y��Hk�4������B�]�0R�}$~|L��  ���~�~����4w�)�Xָ=�Va�!�^^��#���}дG`.ɔ0zlu���ǿ('�m���3m����D���f1�7?t�T� ��i/M Q�ꞝu-h� �Z���\�,��a��M����u�8��i�pt���Xt�ũ�J��5�nA~s�:+�_f��!���l��� �Y�I�\���.�,�z�ɪ�����o��d��;2´"�ߌ%P��{���IlR�!���<k:8���XE����4�~!]�g���5��yd�L%�����-��]��w�{��(g��_2�U�e���E����~t�קaa�}Z��/2����v�W�g�Pńw��x�{X��Tw�{�@�U3_%]���$�j���9���_a���\�UAM��ў�!h�O��1�"�C�g��|=�{/	s%O��/�U���������XŤ=�����.���4�4�VR-���h�%� ��+˜�&��;��^�Wx�L>�e��Q�5<vH�fB,] �����;t�a<���P�R�*��z���C�(^��89���8�(B[�	?�C�zY�o
��=/c�"t�?�t�+[����ɲ���>�2��|��I��r��;N��{(}���|м�0yeC����n�%h7�!�dkLn!�%N�Z�	aL��,���EB��Wmu'䒄�Sx��M]>��g�g�NN����� P��������ꊕ���ԏ��H-�����fろL��E�=΍���p'�i�H�VR�������T��'wsN��7���٧�DA��%�������@Cq"��İ�YQ���� �=ݙ�e[�Ԩ�7]ب(ttQ�nH��LJޟu���Xzf�~@0��.��I?Z�}��ӭ!��Β#B����޵�t	�j��Bt��>�W�����Ԓp6�x�8�Z3����7H�\��c.�&J����,�Qh겳׮�D,v���u�O�$�6�����$z����={v��*��א��	h��$�w�f �t��,��_����ٍp�ٟc�K��L��0vp��T�. N+���m�]�{� ���m�'���q�h^�.:��/F�k�!_9�)"�I���H�J��ϟ_2�:l����o� �/^��^i���;1�j�>�=��6�K�Dr�.$0>m���;�	,6��<2;??�Ț�!���׷�͸�o�����;l������x�����㳝#�\ۏ��S�����^��R��>�L�nj��#ܜ�:�?-h-���)a��v&\���K[ŞJ���O���xɀ%�Z��?���cw�X�|�4��O�4�vh:��EUS
�zϵ����
4�{�X����������� @�S�`�)Ǹh&�z�.�����O��Ӝ`�l�FL���i2�Ny���y��F�21��Z{׌��㨕�Ќ�i��˵�ҙ�".���e��E�(�]\��@��+ ��\�T�RxKk�+�#�dZ�+k�<}���p���%)t�)���P��g|��#���	���ieg���O�+�`&�[k�*)�Vgd�k���w��|~OD�w��5��n����5�OP6 N~#���K�(���3���/R���.k�juI"����8Y��.��C�ss�����ș��2�J��	.�a|��;#B��m����B���dL��u<6�wK�z�yHē�*�&��L�����~o=y͕ܸ������x��~�Z`�Pp�o%��V��%�~8�Нm�[4\h-��kp�*�9���ص60�����闱��G8�aDD %�[���Z���(Ι���s>��y��+�.�����(q˯��oEv��d�]��(w/���{��{>��9�+@��tgK�9mX��ɞ�e��ޟ�/�{�O��|v��q��Y�9��nm�\~�{"���)"���|nO>?<��vz�����*�M�z��X�ޏs�݊�ޠ���@��gy��I8Ԥ�*_Z��Nl��y𜻢��g��Hj�(7C��x���&p�b�M�no�i&�Qi[�g@�/��0+8�qh��dٚ70�~~���p��+]����]�>�,	�\++�Rj���Yߞ�c�4���n�����f�8׶H��������Kw�.gYVWq��<2p��3��^v��K<�����|���C0�{$NZ_���$Tq���{I�@����ڬ���%/��@k��&j0�ss����5h5�ݴ��Ao�͹�ϙbQ�Jt��wF\�b��7��DӅ�!��`�R�fg�m���>��+����a፝��̸d����;�a��K>̅V�����ӣ2MT*�{	Y�����Y	��W���@<�cC���[ݎ��V��w�;���9b��
�E�%i��/��s��i�~oRW3�+�[�ML2�w���{���#̖��д���д=ר� �E��NDu�sV���ϪF�)~�_w��>����nH��>:&I@�$FG�UuC|��!J0���@����GS�o.\�鿨�h�Tij��{��F_���+BA���2��}!��U3��2}���_&�^�.:R��;9���i��L ��=;%e}�n�K*�{�ueŝ��΃e�:�ϕ��ؔi���d{{{U�77��@�'��{�B��ZU��Z��T�*iE����B���{Qt�l�]-L\�R?�a��<?�ɾ�b��s>����~`n�2_���-����y�(ߔ���6I�Ͷ"�i�+.qpH���A�!d�U� 1q�ư����qO`ڛ���B�9�z������N���[���/7�+���иDv�!e� �|�x���+�j��_g�̸z�;���xn6�@W��^�@�Add�a�u�"���2⿸n��!�%�c�0����,�]���^�T�I�T�`֏���)�\��@z싈L��6=�-��H�<wmm]�-�����O���x��֖薨��'XAԻ����-��'�s/��<�dC裹g�g�v��'�
Y22/�ڻ�<=�
��J?7�����w~k%O��77�Y��y�S��ŵ|�{��g��9�WQ1@!���}����"7\\�������CsN�CsJ�w�H�&;@v��J��x �1%dc[l�2��g�Nb�&�!��2�#&t���R���V�'�ÎC��v��� �U��Q�Q�뇱�����}N8�����¨(��?�L��J{��dS����F�^�+XbH5S��R��V�H^bJ�Y��/�a\ŧ�l�A�\�w�	�P��z�O�A,�K1����2���F"H4��.�D!�5r��,'�}X~W�ʜ7�r����ωJv�Ƣã��y&�Q��g���ggA��
 ����I6%v=Bpm$h(�~F��"pc��ɧ����VB�=���y�4R�d&#~�"UX�8�ʃ8a�&�T�ʺ}�</x!ax�,��-���@�YTb9�t���U ���;�����r	�^DIADE:E�KP��[)��V��ne�ai�.�����g����8<��33�}�=��y�O�|��,�k'	���P�T���{f���ec�{�ʏHD��*�/��X\��uH�%���ү^���Yȕ;��G�3��R���j�=sPr�B�]�{泛S����
��<+�$�����^���F���O��4�Ź�&C�\1���с����Ξ�O��m+Xl�����(�:��ڝ�GW���.Pvo��yR��p5'��:b�_Y�@O*p��Du��Nt1��"ՙXP���f�'��p�bvy��EF�D�*����w�?����!Z����!�̽�e5�h�z���&T�]���R��ThLR�9�X 7�����l�����NC/nq�i!�u�O,K�K�+�urf��vk81�ʄO־���#�Q��ږ��9�u�0�X�s�]NW�y���U�p���rIx%�b�	�\�B`� �E��ilS���H��Lޤ]<����h)�kf��?���<�e:@��U�紜���u��:�����7ׇ����.	��?^�r������c�G�۳Y�[��Im	j�c�Mv_���k��iV�HP����v����_�:Z�';�����L��=�C�v,�D�`�����`.�PR�h)+IzY#��p���|ՙ/�1`�bl���՞��rX��<
�xJ���וH�r9�@
�9��Z��-�X��6���i��mP���Ik�D}�]�onu��AU�X���^��S`�{R�n��<�澁��R�7a}���~�+a��k��!�v��1*_�vKn�T��>d7���Tn�}sbA,�%yj��T�!�`sݖ.c��nL2t�w`ʢ/�F��#f8,A����n���=j��z(.��v���:�J�͆rqm�V�� R�;6���他�
��Գ�_�����v�N�\
���$�[��h��";���[V]>?�����1�J�N�?��/G�+��2��`��vw�+*":������w8�y2����zh]'�nWex�Ӂ�s�o��"�-A�%�jC���
]�x:D�2ER��^;�Y%������Y�8)w�ʷ w1=�W�������W7�b��`��Wx�b�vw��_����$�V�*�=H���>dp�3n^ǎ��������xNg֍]Ѩ6,��G=��XM�g�|�@R`�&�#�������*|i��%��P1��P:�0�̧�VC8d}_����%w/o.�}��6�\��"h:X=�_B�6�4#H�b��x֡�!��$�p=S�<�QC�А\��>翻 ��R^�sv�A��{��C����c����R;�����Nj�&̐wpwޙ+���o{�5��$�e��:��qK�9o�8�L�'_rC�|?teJ=1R}[�\�QE�f�7?�j9���V���AJ�ȝ�Ro�T`]��D[�uĖ��Ỹ�����(uv�7�'��-�w[Ìg�*��L��A~�L23#p�����ٛ�:�$!#�Q�t���f>�P�ce���:n�R��uH�Ҩi�M#-�)?�_a���3>��r�.����$�н���3�y��F��$p+]Q:E��	�_��6�^h2Y������B��
�f��S�O=��%�v��T�.�����l,�'������M0�͕n�^�&pX���[ ��
�eʿ�`%���ҥxJ3u�֏���+�R�I\�߆2�bѹqDn�܃G��~����S�p��#���jSH��>N .T��+������~��?�U���Zæ�X��HI"`-�?ɐ��XHov��i�"���AoT����UЩĬcUSw�+Y ��q���eN�� )E2R{���ϟ���gu�_��\h~�(��(n/<�:��Q}����� oԕ���^iW�_���)��S���=�>A SR��ʼO�r�0�?���+ʚ��ߺJ��n7�oq <+PU�P�,cN%b,�*��\�8��ܜ!_��l�µ������<��;�l�����c��_���V��y:�$�^�ٟ���`�(?�n����9>9��6����k@A�SjkJKk��\�MsYX&c �&�+�Rb3S����ŭ�}W@�g����R�#�����	4��87��W�8�i�"�.�ꁇ���V�����-U�>XP���/)9c��x���U�:��r/�>�}ZU�v����h�Z���a`��Z��Y卺���c�W����acK��Xp����6�Ԕ����n�H��U�',>��7�nni�i7s)�ھ=pK�Ǯ�x�wdm��~v�}j@y�����cƨ���NsC�껼�D0�sڕ�V���}��b�)�[�L�])�FH2�w����2MȪ��>|W�� h)�h�?ɬ�c�
K׿	S�G�bAA�4�@Vf��.s�^��w��C=O�<t.M����9�-��fG##E�����V��V��-zn5f����MZeE���d������X�]���l�H�+�$|q+�Y�!oS5�GE�yr��x����G�kD/����M��yv{j�uu}�;�&e}R㒦���lf��=\{�g;U2����M*�.ì-�_�%#����u/N���6ܘ��!�	`=��>���?�(rm�j=g� |o�
sq��\@ѨUځ�1|7�����O�]�bN�?�Z���,�T�$a+JQ��{D�Sw�b{Np�D[be������^<�ff�}^wE�_!2�$JKH>V.<���݁�'����� ���0WP<�xo��U�9V�l !��j�VE�����	�:�~JV���a���8s��_�|�tg~f�1%�.�θ\<f��r��B�#�_�`_���*��7F�#JJ"�"?IJ�&��zIAu�Vz`����yHXϔ[�A��ʕ�=���K���hA�"�2$����mO��]V��[�y,����~1Xvp��ZJO���P�I�j�?՛���~���qh0�]�vv�=7u���j��=�T��{:UfffeT}_]�:�HV����:�d��t�>���\A��I��	�xn�6��{��>I:Ï/��i��h��!�����6�#��w!_���8ި��,E��:��'n���
��k��-�3��9%�AJ^��,--��x9�i�1DcՐJ9Y�g�6���콳p����My"����p��v����ڵ�]�R'�E�s�у�3�jχd�/�ʒ	!�㉝jz5$İ��j��E}֟�󊮲3Q�k~�]6X��1�������lyg^hE`vN	�K,S(5�&Z`��p��k�����,Ht�颣��	�%�A�n�ey�\R�����s[��d�7M$/�9���qN��r�}������T�6������5��L��R����&`$�e��GP����И�:�kH�W�v���W���\�°�ܯ��q8-<e�_�"���ú�~_�������ڠ%����S���K������N�����n �������:_1��*�t�_�O��˟a�myn7�\|��@�$ �	
���4��9�Y�������acl�z闱��BC{�):z�_��Z\����șt���W��y�ya� t����#�|���R�4�]�҇^�O��g�ӽ^��`��"�AqK�U�T�຦��M�&��jF��c�}�6�g��u�~{C�'!!�b��?��� S\Hn ���K��]AFy�O{O��13��/x�~y�- d��+��<N�e�O2!Jܕ0�s��S����8�?���W�������~<��n����9c �4�J���q����p�)}���oyi�.�;b6p<���Og�9Z�O	B���>��֓3Ǳ	�
��|{�x�.���J�	��|�>=zqUf�Di��s������y������P�����Bd��nD([��x�)��γsx�R�*����BՍuT�\�^$�O}��"J�0 ��,x*Ͱ�������m������/�MG����cy�M[��J�Q.{+�-t��/ar�[����V+��"��L�e[2��h��
cVr���TY0�D=��Q�3ߚ����M��P�{�:l\ 7u$�V�����~70��Gs�W4o=qj���y����7����f�����1b��D���XTbd�T˩��Y0�[\��tB����C/�`��)�_�'0��d1%���I� �y�|��ı�EX�,�+��H�vu�=�7�rƑ�ii��y9Q5N�s���:�v�L�n ��7����4�f��(CƧ����v��i?�#�����Iۅ[(��9^[�_<� �{p��2�v�d�{��|�)�)����1��$Q�2rEV����@�C^G˷,\��]y(��m�����,�Wb�����w��ff^C�C�Fs�2d�F�
^$�\�++�Zδ<2@]����\2��0��¨+�Pj����F#4������*�ǃT���P1M5��>��eQwF#�]�P`��w0\�̬�&Es �O�������.��*j[p����������D�l�l5���R������4�D�ܲ�Ng�t`����/����<����ꥊ��;,D��������!J>�4����}�s�r�����l�;o2�MM�JA�ƉWe>O�H����-�1]���j�k�[3�ƽOGmq�#օ�2��+����ػ��СV�d"�������$O��@���V9�0 ;B�11	�f����ZWG��LE`a)��1�(}|܇����C��o�뫬���Q�p�/X� )��n�\�(Ri��:�=����f�~-�	�[j�Se�$��{WY�����ʻ�������z�v��`e���m7ƿڵ�.vx=�1L�r��@����vK�z$c!]*\�ݸ�j���щ."�ә�%�d�EQ�c���\n�W���j7$0�'$�~r�E�N**E����?aT?{�ۖ�,=ѝ+���ji���]?'������L���~��m�e0�����:�������� ͆����}'!]%:rM@�8j?R>����m$��~��4T�`�f����촄_�Y&�jj0�r�s��)UB�'5UKk>��iT/Z��>��1G�%Zq������!7~Y*dr�v<�%�	��O�wR�6�}��t,3��H��ٵ��УNH�zc�1��~�-30��[K����D�K�Y����c�)�Ƴ��iN�t\�&��B��K:(��������M�|,�_��3MDw?WK?�r>	�l�[�|h3mtL���v7�rѱ��0J�'7�hՌ���yd��2��[�}��*>���?Cg�Fg��{	
��Xo�#"��AR<�/7W*������j��� �3�)�~j�<X����)st��}��?O��N�Q{���`pi"����@M���/���آ��r+y�� �'n88��8������{tq�Q�L��`@�q��w>vf1wµSR������i�́��^����+1 !����U�k2J�V��� ����F�
�Ry�;Y�O11��v�_p%̿��*b\�;��A2KlSIme��6�������V�"�����+6��u�ȫ�Ulum0�'ǽ"��SS�~��)�r1�U�K~qd�˺���i��P=;Zp�x'&
~u�n���&|�
����QYw��7?�bLZ�[���Z��k�U���ANU���7?uV�t�?׾�؛�\U��£�Bub0}5������{Չ17W#�$��ibl�(���h7���1+�ۈ Z������c���?0�;!��6<�uu� ���Ɛ�GH����&��B�1ܟ�S���|�i˪v�x��6����	��dn軉sS��0�N�}�ÅI�,�,���b����i�!���� =�l�g
`�|ߋ���'���N+=ۋ�%�M�0(�M8m��4+�g�!%���N����i)7��Bk�h�W�n7�����jq�����+$�1��hL�����K}� �eU�!�Rp��6i(h����_��s��
t"2(J��������C�z��Ps�߰+}�wAJ'h16v<�n��Qا+�2�b��s����_���?sD�$dO���M�ڝ1����b�R�s�ׇ�%�.³Aj���W����X���V�7���#��]ó�h1팒s���x��W�\��8���pMM�ט�@ʄ���'��F��!��=X�@W#�\*�[z�iC��{��4�I���?b:�w�/n�!eE9��{����3����E�b�H��`-�+[^��Aly���չ�Fͱ�>�YJ-���(��F%��/:�dp��>�/ ��x+C�^i	���q]I"�9�B@?,�b�{����Xl���h���B���i�;b&����Y�J(+t�!����Q��J�Lzv%����Q��F ��]���$;(BO�Ř�q���yJ���FY~ ��T��s6�â��o�i7�f@~<[���c�>fwu�5��`�
��7�$���%;32*��DCuL^Du!Q�y�C*��W����P�E$����W[@�H�G(o��~����������	L���P0��b`��tH���]NG*ͨ)�^ڌ�����jH�A��z^�xu��&�aK������#�Q���Kx(�	k���x�u���T]'�v=��Z��=�DH2�����ю!��\6�}�Y��gDM��,�5^_w儾���d*�ۡ71��[���F�+��>��2��1z�V�.�'�t�2���,YԵ��BT�ʾ���f�?;Y]�^�-6]��p�'��Ƶ*8}T�����݄ZqSdi'N� Fql�i^��::Fʑ�}��t�{w����եW-�������nNz����G׀Y�,/+�n��e4�!?�eB]���Gi��4-��e�����3�~}�!��R����MM˂Yh�δOmIr�����-'1��
'��>��9�n��$nnjcMҿ�,�1:�
E�Ʀ�g���)r�\�����ec�j��n
((*�]���ϳ����G���9��,/�����j�t�j�rt������ͬ!�؊P��6�`G�gᣓ�P��Ĵ�y�'A��G(uqޖ���V��%9�2]�=��k��bu�5A�{H�]gwp������7�!#Tw�m;]<�� #D�Y�tB`J�6y�ܟx*.frd�Re���j֑޼6�]1}��3b��C��(/��ܼ�i���>їH�|$��yfq|�'��M�.��,�_fNM���?"$6R}
��9.��@\��=?����2�Fs;Pmj�023H�tv��`�}�������=���Ѽ�#�d��
2��ݾǏ�����?�M��s�!��bFjB�\��O�J�r�񣝣	�TDLfU	 R�r;I	]��t��F����_��n43#pp���<ݛ��BÅ���s�0	�\h�����~�L�LKН�^9y���'�gw���O�6� ��P�=��!Y���
t��9 #�}��s6G-�硰(&^ݫ|��{�sQ;�??�iv��귯��jT�{�����d�ٴ� 3������*�,������)C��kdEG��2$0:Y��\Kh}�a�3���5e�u<\�}�-�#%��)�1���M���Ѩ)ٛ%��"�Aj�~�0����۾�K�ٺ FH!}�`T�����T���L�9�G��|㪛��Bc��EF���|�I�\9����Go'O/;?u�7��>�#����� �D�������"G�B\X��:UK�����DU���_G�n5 �%��SqJ9�tb_ϙ?�����j���u�yX���gCE���M�:�;ɫK҆�ӹp�`��Ų�.��zL�? `�E��~�]���}�g��L7�i���JO'V�ȟ�-�L��h$rKCS��2kԡ�=d0���A����ht�J3j�~<��}�^Q��6�РP��yy����du:��BQ�">q�c%��Sn�t3�n
�@����Ё�z�T�""G
���dyu��I�:�Zna��c�a�b��I�2R�g�Ǩb��\\�ڳ���kS+�1٣���(��.�H����b�v����>u��ϝf���7Ǥ�p�<�BG!���M<�vO��NIɰ<mi��8����}�������W>�u��#3k!��3
�MZ�΀����8���<�a�Td��r 쭿uBr�!��奬�X�m����&�z�����&j�8����A����Ŗ���ezŬZ�}J�twG)����D���ҐŲ� �u+������̼������w%��| �b�	2<s:��D e���p
��5eܘ����!Jƕ�w���͗�>�U@��o��/4A�o2n�|y���P�6����0�z�����8�EeQx�P<1��~����[�g��b����a9�$j�n�ru-��=y��=��5Zu!�	7ξ�7�i��c���!DI�2�X�K�!�][s��w9ZT�(�ى�|�N#"/�2@�a�����P�Ú�Q+��it8Q��;R�#WN��Z�'�)� �	��B^M��O�vg�nIJ�h�Ҏ��#�	�7�]��?�q˚��q�5�!::��I��%srl}�����5h��0h���"���us@�*]"J�si�n��n�oM����u`
Sj'���f�~��h�q+��i�ٹ��l<�X,G�����u=��Jz��1���p��Rɏe#r�f��6��C���I�de=�v�2��U�E�������8�>�@0�-�b4Szo����Z���M0���_�Y4���ai47/M��T�cb���{o��#��D��guL�rۉ�YBDީ E�!P!'.�O�u�^�XLy*`x{R���?:��ۼ��7���1)RP��|(J_��Д[�kux�����tEEE���c@�<>�V2�+H��r����S�����ǒ�W�>�	_v3����+s�Ю�ANŝ眸a�)p*��H.v ���1�I���En�3�
�I������Oo�b�t�u<��\rW����0��V&����pd���[�ۨ��eSa��I��mU|�N7��!D��S��D�ff�,|]:P-� �ws�CR��lT���M��p���u���}��U��ڋ���3��D�������bP09M'Q�V�`�.~͆��'ׅ���B���^�U��(�8�}�3/�n�ʿ�!_Y��:����P�<��W�^��z����7�4���p�GU����	uvu�H=�H=��zbS���$ڶ�:7�é�Ԭ���آ�_�=���1n0ra��d4��z��F�"!.h�I�Χ������6�F݉�.vZ��<-B�{��'�Į���&;0��YoX��n��){��Jt���g�H;�W��@m�<m�R=8OS[�\Z�ȵ�,��j�g�c�O)�1ZS%7�+�>Q�˂p���ӳfoH����AA�xL�<,�m���.�B^�i��1ϒs��kOy�<�!._~8-����-gv���=u=L�~{i)�q)��F�����gVK��K~w�ܷӥ�-3������7�R���E~@~��g�y��N۾���B���<b6��,"�bk�'�C3�B�AY:>�#��w�Q�و�P�B�_4��qX?c7ư�)o��U|���|	��o���V�Z2�h<�?���U�D��o�va��?y�7P��_����W�x�^���q�װ� �:�֬��u��Nb&D��|�%�]�r�oENR9;��ȏ��߹�8�������1�,���	�{�oLy��|���Eb�Ϋn��%f'Sm�*O~_%���^DYu��Xy�)XHz���Aj~�(�h�q����~����0�v����2<xx|T���,!��)1�g�w\�L�G_G��`"`��[���*��h<"l�2j��pГ"=nNBt��>���SX>ɘQ.�U��HR������ގ�l���M��n����uԄ�b�� d�z��Sox�[~p=��*�0��z g��K�����/Ưr֐�_��a��_�)B	�-|�tq���i�����W��Xd[�Gw?���6*h�z��x4�(�݉g[���=duGr*U�?V�6>6�L�ݒ�����_ۣa���	X��n����V�̊R��l�5�+.c⿜6@�����ƙ��;��yC�^�-x��VC��WI�n˹��5%�\8E�V�?K=.��埏��>���$�� �ԛ������r�o�u[q5����O?���DM~�8�۴���=Q�,�u�$�{��H�i�:�9�����Tkn+�B�D:S��ϖ�ͺ�5
z>�W�E|���^�H�VK���1VFRϛQ]�*���-C�PX�^s�����B�t���iːV���;7^�6Dbt����/����#�Z*)b(�(�!H&nn.P��w�×�x����xSS�`�%�RS���I��P��оJ;���2��c�������E�+-���P֨��0�e�1�r��̮�^q��Œ{���_^���\;o�5����4�
rΈD�^<�j�V���[`�����җ鍍|u�t(�P���C�$g��q�k�qQ�)�`���G[��[��B�M^�Pp�DFy�{�����>�0�E������z�gޯL\���2�V˪���x���NK����S EQq����$�[<[X�m��tk�a6j,G�����S���b9Y\Ћ&�:��;kW�d5�;}��#%��,M��mr���11C����7[�/X/w���G���O��]�u�GX���W��:땓%��-��;9O�yAZ��#ڠ�@���8 ���q����Q�rλ�O8��Ū�v�+�2'�&u�pQ?�2]G�4%�*���>u_h�a�k��p�Ͱng,�5Lo>��x���ShS����;�D�l%�؉g�)o"��*횳G;��_cM٦qJ��mp;�	A����}KLO�m/�����3�*79�
�jN�q�e����e���mw��	 ��ef϶����p�׬wd-��C�����Nl<�Ȥ[����� �"N��	.G�pt��%şf���)H��ĸ�"7W`Q -�C.vH����q@]�x�jd�!��� s��9Z��F�پ�Q;Q�W�Q�̋���3h�5XcY�`ڝ�MA���Dc��dl�^���*����"�A;���iFT�G����N�]Y��)�Q9,�4�����4>�y��g�on�vN\��C2sN���"��$����������J�j&Hm+7�L(I\)_t�}(Ğ�Xf��T��j�UW�o�9��S������GGY��r�ŝK�5c+G���'-�J��J^���}�J�i��Li��!K6.�����T@Hb�#�K-�)�~68(s����6B�F˼�UJ.s�V��[�Y�B�N9Yd|���<��Ȭ�#F��{���qv ����"�dGs�0���>���i	'.xo75���aA�ؠ������v{�岽I���M�%7��iT�9�}�snX�h�7(���ѵꝦ�	ӿ��{$cŔˋ���r�����I�U!�mc�
�G��A,�?zR�/_����@�#z�^e�."�n��i:LG�����A�a�����\�{+'���?��nZo��VI��9Y,B7���@EG���v@P?"��Ŵz`��J#�T@��~-WįE�H�9����F�m��Z�R�����J7^����;"r��A���.R�@	�C�1ж����mm�\X�g΁��,q���-»\��/M�
�F�����9i���$���x��ML�(<�k�dC[n^6�Y�~���t���9CT�T��:�V6҆&(mdt� ���m���!�G���4�%8�� ��̓�?�V/+6����Z	�o����w;�[;ItݖB��aPQV�-AI���� �����n5�s>�^9��.��5��@+�,�L���Ifo�b�j��ˌ���+�����OI��;Vbb�]�q����K:&S��Ϲ;0u��3��-d%}��E���� � ʶ�yq�'#)�f4���  ��θ���,�����֋�P'��Q�v���"��KpqB#e���14T����̴��#�5��*�Pv�����i��a�a� ��gb�
�\��S�o�1���� ���w���m�iv�Y$K��&-�;b�</��fВ�R�d�p���o�o�b��E�>r��4PY�L�#�g����S�z�?{X8^��B�[�Q4��TZ    �֕�7�������G9!(�(���ZP��G�a�+^����r੿6�9�O��V���n�
��K����dBU>*���s���9Y|��!�)|4�AbΒ�1���j����w1�7��r�-pO,��7�+���ȣ��[	@��'o����fB�ŕ��x�I,��� �u�nA����DS�`%P�
9���x��d��ø*s��.���V���YɃ�)�E���{�E�JY���*�||'��N��R����"�;��YG�l<�Rt��mHS9g�^�,�a��b`���=\���ѯ�tB�w�O��Khh��~L��uy���� �,ʉ�JYq��
�y��m_�~��v�]OĎ��������� h���娼�ҁ��J�6�
�(��&����`*��<ˏ���LJ�-���{8�h����i�T��M�9�F/����Ncz�k&�b� 1I����y ki,-�p������x��L�@_xT�<���>�pM#rif��m�,�lǂ�����~���:.�YϺ#�� ���]kF𣰐�**��Q�Z��vʼ���u�D����^��n�����b�y�d���M�l�Ҩ^-�w�e�(�x~���pg���Y�G�8[3_���]��`���Nօ�>L��Hgݮ�p��Ąہ-����әRͮ��T�p� 2�:��P�Q�/3���~T�߰��^E#����<��@h�dQ�ו����	|uhzx��<��r�w?K���'O�Δ;w���~��!G�����uU0���?m,���(,?Q[
dܷ���qӖ nTt�<?�$о?V���(��P]9{}ܬ������נ���N�.�\Ov���Ǿs3\��ڸ�~ �iA�1�G����X�I��&��A�m�ϡ��-��Lq%�i�+��3e=NFI�*V�Y�7�O<9"�ac���1�L�)w�M^&�.eX �Дկ����j�����DD�SO`D5������%`��Q�j�I?����`�$��`�� �n�wet�����(��K[7<���n_11��!�%}��b3�PGqӏM�[h?�ɐU�[����b�15^\�u0J�U�V�����}�yA���	�K
Uj�>W�;K� U�܆�-�'�x%@׉HOײ�U�8��jm�8�[gLdt�h9='!���]!�P��]U6��H��j�f+�JLǛV���U��8�:�1�M�4%t��%t-<�;m�t��h*�|��=(�K�'���i*Aǌ�8�EF�;��� �8܀%�&�Wr�L~~�V!��R�B%2Q/r��dnC�k@�U�RwWב�󍍘`�sT����Q�o��,�����\��w�,&Q��Ѷ��Ƹ��&6B91����P���<t�y^���uT'����0���4��p��i���`Z̔9 \V��9Pԯ���6޴T�<ݖ'l��$��d��2��RS.��E�1��)B�7�#캊�7/`]~ ;A�Y� v	��Dpo�����*Ɔ�8g�����M��n?r?��,A}!MTaM�h�MEN5E�*��<���hV���.���婤�蓒
��?�+��1m���N���h|*W�Vjl��ԝ��;�@�/$D�F��%��=��)�I[PR��!!��66�>��;�MB����o�Pw�4>^�ML�ء`E�����v��ˑ���x�n��Z��8��혤Z����m7�=_��p�׻��{��iۣS&��%0����Z��c��){�-:��D�@�a��^��	]!���3-�6!xO#��7�.8O�Wn�eVH��j+	A%e�~� �b;Y�J�
��a!
�GǕR�������#L�y��q�`���N�~�')�� <+����_7sd��Ɍ8��� ����Ӧ%� �復�zV`qf?n�M9&H��j\H�B��MUC�5bl���eծSS�v�UӃ�^�-��nωUx��k�N���^6�UT�T���u�
h��x��ǃ��.�>$�yV� �0�_�ʷ��̧}�4O���D9Q�va�>Ww>:Pр6���O�n#�hq�Q�>�׊��jV�@آQ�Ɂ6ѫ��b�����'(rNǯ����]:AP�Ol�ٚ��h��!Ѫ��:L�P.S�I:�O-Nt��-a#5��!��M@�N;#-��=��P�O���#�ӌ
_�ĸ���#�O�n�X���;GXnj55��8����~��U���^?w����B��w��	�л�� ����Q�Z�'n{ykG"�f�k��Ō]�R����vp<̂�=��=ᆛX��/�X~�L7Y�}e�c��ƈ"��
v�5K��ը*�q:ݒ_H5/�h�(�98,�����
`�ffIHjoy"E��<=O��s{�R��H���vff.\�����ꏖ��_�^���a���0\Z�R�7�"p��Ӄ��y��-���I&T���<}@Vs����n�[��c�C@�h���Dv�=q?[q@���PVn�p�,�V=�'x����x�۠������9���V�����9�'�Ϲ���Cm�ﾜ0gq !���[��kk?D��(@�·V�D���������_r;���%�"	�I�D�ftT푪��kh���5V���-�vz��R[ʏf�29 ���G�P-�=�'g�&������2�Dk�O62V�$o��3d��O���4�߮�h5��U��dz�;Ob��g�
0�F&�Gp�	�r��Be��"���m�
�67'���':�-��;�?�D;������5XOԶ=��Y�F�^�tE���������À����h����7�٠Ɏ���Ɇz����2�(m17����C�n���[.w&1�k�f�Mh�.X�f���1ݿ��eh�Ȇ1�jn{o�e_�Pff�����6*BK'y=�97�%pO��HV?�m���A�����S�bo��{��Y=���aݝ�"V�������E�EdJJ���JS'w�_{\�?�S��K�c@�YO�RG����N�"���2�+��%���������nO��*��0�Q8n#ë����}d����@��N�TI���߀՛�&]�d#�@�9:E\�J<�k��P�r���SV)l?�t�J�����i�`#��^g窜�d���s,1gϸ�����wn��(�Q	֑-�tq��B���`ny;	�����G�kif#�A�������|�v��Y<qόi��hW�d�����n9�����T�ҥ�����c?Rz�VJ��C��:�Z:*�8�>p�h������������:Z����Y�9/y�qt}N��#)\�I���sA��+C���M�/��1�8��ݜ:����8� ���KCh{��.	��mN�ڿ�ԓȫ�r �JK:R�g�&�E�J����jg��	����n��|<;�V�M�j��ng���@_H�huc�)�Ӷ�\���OZJL-{g'$ViS�u��s��[���(qH�~��a/�BQ�$a�m�2���?�T��4��~j�B*�N�w�� ��|��OB44�TW�W���FrwӀ�z�`��=�G���vT��{�m��X�Y�v ��������E���0��1�`\����ЕA�ٿ���Y�sw���ym���I;x�c9�&�(���z8�g�_��=�2��o�
mJ���P��/c�o�gM���?��������[j��ں�J�S��i�aRTp��$��(�d�U}�ͱ�i�M�٪$H� :M/��9YO��MOM!EV+��>W4э�늛:;)�.����^�����#��z�2�����i��}�����F՞f�2�6<|�I�FJ�E0D�]q]����o��Y/ʁ�EU�6�"GZ�F:�C�e���_����ڭ���2�+b0/��t@���E��'JF~�����(�>��5���a�Ձ����ۀ��r�!C�w�����Do>���B�Ѿ�v�T�S�]荷K���$��D{B��x��UGG�rSu=ozb��������3?��*�9qvؗ�Ϭ�� �`h-o����Y@����d�
w5�B#�;���PPgS�ө7��?�r�r{d�[��,��Yq�����9k�C_�#8�3
�裣���Y8\u�p�9B\��{���}SS�B��(S+��ՄAդ�Rn^�\^Q!`�����y�%`o��Ȁ��H��<_��z�j�!����R�� ��8EޫJK�}���{��v{�_������H�F-����l���5,`nn�d�G�/iU�_YS��f�n|	�G��rҿ�^T�'�z��4��U��L-rh/���R��ɉۣ5�5�9!@2�w9 �c�e�Σ[�b&ȹ����˝��3�s/��#��?f��������r���j��y�HL귒E�[0����e���K����e,T{F��H����Clz:�Y:�'}A�L��\���ѷ�>t�P'�������xyaGiE0=��97 �z>R��{�V����1v[��CDŅY�j�$��Y��q�`���2྘����	�k��@G�ch�ur��0a=P���%�a���o��<�r���60�uKb""��g2"������|ǃ���\�DK��N���7�@IU�1��A�r�w��E}Q����C�:�_��n{�v`��kJµv:O[3wmD1���u��F���s��d��g�?��t�]���$i�z��*0 A�<f��_u�Iw��+M*���3��*�KF}�ſK;�Gr:���h:'A祬�lH?/;�.W�.����c�nC��C����K#&�e�`e�2x�᭭$�����^����G� ��j�9�}D�,�M����P�"���"9@�T�O�Z�r2g	�����BET��ɮ����9�A����
��R֨��rҧ���-��o�im}IB�ݷa����S�d|N�U�d��F}�J���
��g��qڬ&��3= u� ���d�0Q[+��W!��2Ն����F����0eӂOrkf�ڱM����7*���xLi?$d�g8+���,��+���-��Q6�ͺ-�����I�ˏ݄ޗ��v�V�	.o������ݐ"`,Ks�$���Vƍc�` �́�c6Z��TbteU����5�޴��c���N�m۫<xv�qa	q�g�1܅���������2�uع0t�d��{9d��FI�p���t��0��u}7j�nS�<�M��������7�R�T���b7��ka�ग��ww�rV^Q�`�:�N�Œ܏�Ry��n:�y�+����FDཱྀ����x��R;��b�۵��e���ߢD%գ�;~~���0c��5,�f>�����I��p�����̇�`u:TN�BB�����P*͌���5��������mZ�8��V�d8�aC_s��`z�������eIvܰ���R�qF�Js���j�VHJ�+��jಉ{�5.΅��g�/T�0��H9��.����;��<�����04+"�T�l�+H���t��1�(E��t� M�
H����A��������K�<1yvޙ{��;3��)�C�%��<E�e#'�8���8aR�%��p�&��rF+:n ��u2�תk��z�<Y8G�zEEm׉�;1��(�9)��i���X����G���=E"�\��]�UK�'�l��.޴�7(��9�88XCB"��k�s�K��Y�i���<*Y.m��C�� �x"y0}���Z����Pob�{K��{J
���p���#t9�@b5g�Ͳ��7$��%��r�~���<�II1,�8 "F�#��ĭ�<O�hm�w����\Ά2쭞��sl	���A /�.����S-Ʊ�yĚp��o���x�F��FZ>�e#�(�N���D��@A�2^��%6�oLbk��W15�]@76��)�����ߛ`�}�8I�{waJEzv�KM\X��y8�PSC�|�����������"��{�ap�M!Rh{}��cK�*zyܯ`��`�6l�=��h����V���O��4T�KW��S[Uz�}0���Z�Ͷ��F��\����g���Ȉ��9O�S�V;���BMήG�Y͗
�b\�����B�l��)���.e���	�d�~0���W�+����?�c�]��f�>4�u".��l��/����D��Esө�c��BY{|�n� ~I���V��N�nQY��6M&&�����C�~��8��i��Z���Ы36�t7�tnY@5����m
<���F_4�w\�捖t zN� ԕ%���{x�ۦF������Fb�M�� �<�=�%v�KRH�v����$K0��P����|5: ����	�"Jn�}�ίB�Vo�%�D�FF4�͓&;��c��b�a���v�${�$�X�g��E$���� �Vz�������_�NQ�����ݜ�W&����eNY���Ձ��ӺD�C��($c(A���e���3*��Rw��W��;!��b��2-ҷa�4{�xX%�$����Z�Dj�f~����V���䎼�~��|�R�����+x꠼�J���%��CM��~|۲�5O���๞�����ɹ�8�7�w�V�6�9ρP��уM���cK*@b�\�޶i�FX���������e!h��G��g �а���΋�~����\�t�wYF?2]�n �Cw�� ������Nܡ�BAT��è��1i��k?��B�4�`[��W�S�VX��ş?�DϽ2޽��w�����%��|,2j���w�7A�4���S�.���i0q@�忴��ʋ3����n�������U~�y��rR�?�u�<��tK86�\́�� �ŠF�qG�/�q���Iڻ�Ѫ������b�pY
�i���,MH�����X�Ngv�::8�Ļ>�h#Z�c(`Svt�ԥ��͗rv �Y9����1�-:6�+�Ӝ�֢�Uz?����0ޟ��Y2�K/�;.�=&�.JJ�Q+�#���r��hW�:*\ĉP���nu|R��=��=�cc���o�'�J�?w!{o��H�YG`U���R����镏?�����;̨���g���z�6B�6t�3$��A��H���zA3 �9O�C�.��ď�њ����ƭ�p���}�^�w�ѣ��	7���~�Ue��BM�:�7q�8�M_P�C�(���z��_1�� �˾�����'G'wCf3ʤ�F:Kڒ�E�![�����әz����W��Jf�أl4ZAbS�4m��)�[����/~{m�,t1԰��DD,��� U��7lGߊI�Ӳ��~�	$�ݸ�b����B�L�q���É�)�$W<}�i�����	�������"�b�g,��Jk˝�A�"�BBaP���q��~�x�4ָl�������Uh��SK�N+�<�m�r�P:,���J��ԫ������O�o��DD�c��Z�g)ҍ�I��޾�I��g�n�l��r{zvFYY#D4��l�ф�k�%cÊ�S�XB���%�n��DKn/�I_9
�+Nc�i��79�v}�bB�ϲ�l��m��`x;hy����T(��~�$�c1��Wc���S<W7;&�s΁Mk�Ub�L}7NL0�	��(}\nQЅ=�LK�$ߌ����c���,�\Jܖꇬҿ/�EF}�q9���i[93[�~�mj:�{PԱ�d'7v�
O��1}�TDa���HQ��F3xz�kwg�����&�R5y���$%Y��D��(����R���y�E���뫿�.�hu���Yƈh���c4����Z�����߅�� Q�,�8�hП��� ,r�5~{�:!�-�����}�+��K﷋����GY��E�{�,�P�r�Z�µv�ŋ��ب�^|k�����!���{B�r�7~��a6 �}u��Wbj���2'��vᑟ���i#����ST�X�"b���~Sîo�tC��X�������jf}�lM��a�E_p4Ɇ���y��Ҵ?�N(Ei��U��B_Q�Oo��5�.0?��W236P9�C>�x���.�_�ca�Eu�67�i����Q�xz슼:�|�v�7�_��
�Ѷ�[�|��xVԞ;��^H�w���C���Ӿ6e1[m�0�g�s�P���M��4�1���`���ˁ{��l�ҋ	� �� vP^��	��aߠA��K��}���8�8�Gܹ$�^rcB��2�N�� f�u���%h>���EW�a�i׋4p����Y�G��^�Ǯf-�T��������}y=�,�*eVQҟ`ө���q�$���q�w����@�����Bm�
�l]����d�%n����s�COA�����8Q����x�=<�u�����\'��.�	�JI���z�$�t4�5Q�_p��!�=K�|���W=v�K�±� ��cg!�]�~��AA�����B���6�y�V���w8(�Z(��V6�额v��ފϵK���K�Y�|�1Rػ��ߎP��r��&��P��<����갈E��[�t�wD����I�;�jF���yc/Q��`+K+2�h��\
��.���r�:�`��Zb�X���ŚTib��xgB
`�v[VA+t����]������@��$*��ǆ� ��#��.��.��準}�M�!hEޒL�3"q[�v���e�G?�D��on4A��V2�(�qlY�c�(��H�L�,��]\�֬���i��¤z������4ɫ5T�&��wYD���:�z��O�W�l��>�P���W���w�S�I�NPV�����p�)tDu%+��!�}�F���l����9����:�C_�p���Z����z.��n�J+c��ӈ����K���y�h��
�'6�}g����@f��������=9�K�Iv'�$L��e������]�s��SB�y��v�E\�7�B��wJ�}b���E$�4"i鸳�O�r�������Ob�:P�����B��v:��K�	��@��7�=>�m(�&�a���6@E�r�E�c`��U��������E�ӯ��h�B�ÍEZIc��RwG�s�S�En���$]�tjrD�n��Ŷ����=cά U_tɌ���&@�b88  q���Y�F08���1�[ �x|����x�;�-qb���'���us�Sn����q܉u�n�!dkϰq�~��e@�hlh���Ǣ_�l�!:�㝇�����K�8%o�x
@�����}~nl�!��L���'
���5x�����|a{SY��2��gP���x	vdа�	w��#�IJ������ P�`	�-ЗM�|�����	�|�އ�a�e���u����c/V�b�ޙ)v=X����s�oEm�6���H��]���aUA�	��l@V�h��o�$�l�/���^_�����b�+�;��aE�oT�B��zI�<7N��йW���.��Ad��V�i���ǋ�	2mHY3��g�+Z������
�3�,�;��I�d��N�L�b��j{��
�y�ڤ�^w""6b�������;=�e짤Y����*gAڙ/���9��J�d�
�ׇ��7{b�ݺ��,m�1�Qo�8��3$��g}5?�H���WRc�G�ñ�i�{�(�-�[��������o�h�q�����[F)��H�[����|�p�������E]�^f8���+t���M���,9�H�[�0���twgĝH��-F�j{"�w��B������1��� '��I�c��(��;eq\��zn슈�d߾�~�;߃?�z�J�=I�'�I�[u����F�XП�9��\Bͩ���g�T�ywR:���\t�K|}����j�7���[i_�/ǿ9_^��~��(U�߳�,ӉKK�Gq0���b]�~�u����:��k�]9#��P��Y�������W��}T��y�:)K�rDq����܊�I�pɩ)C��/�6�N��a����5��m���}�����(K��ݑ1H�1�����1���(Ov��f�!{��N'zZZ�o�^��l��N~�f�:�%�V���B��VL�J.瞇Ǜ��vvq�g*��abd�	"�����������/0)c�����Nn� �8��muu���J��׆�U��h}��W~׍�.;�z)���\����\�f^��4�;{C����;�X�C��xx��g���k�՚[+��{�k�n�̺!V6�T`��n�f����;�\��.��Ǝ9��^֙�n�*��h���k�:��Yп`=g�Mu?��I2�d9,'�z���/���3H�����#�Ǚ��E%( 
�ru�s�%6v4OsZ�/g���۳5��s+���[�Lj�}�kS,��dh?���&Ox��;�I�����ۛ����[[z����AR&t�_ъ7ܰ�H����/�t��%f��l����Y �/`E��9�}�DO����
�s�4�W��g"+���;�j��>p��
6���ٕ()��~��m��{E̋��y˓����V=�է�O HF>t��k7VBkC����|��lt$: �����⢞5=�^o��3��s�Sw����hh�Q��`D�~����C%R�O�I��SzI����/�wϊ�UQ=�?��c'+�$1�U]=����,��ie��L�E�E6g�To���4�ܲN+��%g���f�x���jT��-!��ِ�	a��C@b�m]~��4d���؝���[�f�㑕�X����>���a�m�S�Z�f惆��U�"8/8��s�	m�<���j�}���W/��m*z�.���{t��H�-A%;vT>��JxR2��;`�귳	ņ�ev�~�	�q~_���oB����Q�3�x��c���'���*]���#��s��I=��e��\�H��z�t�D�{`��qq5!���ƛ��[[�7���}1�ЦT_qZ�d�![ ���!:�F:�M=
�r�D���ya��{����b>p֤dۑl��#�
�K.����=f��*˗"l��j��LG�:Q(�V4��^i�S��s���j�
 <��rH|�r�y�
S��9�)G7��[I�81.���\�r���'��tXa�23��c���dLA��s ��@����_������X��P��CF������b�B��)�az�J"���ޮ]#�{�����)�Jzazz�;ү���1����e6zU���b����i�&��ГD ��I���,	�.$�=�-���tR��q��{=qU,H?|�1buu��S#�T�;����R1L���g���]�Nv �Z��]���;3P�.]:�>1��nn��Y�Ei�fxlF�������glc���:2`����hii9mp����?.FŒ�O�f�LHg�L���Q��<�J@��T�\���V�(��q��������8�
Б'n-��e�@��<�ttTQ<�~un�� ��\��f�O��.;�0 �^��YR��[/����BE��@>(�����!?�ʙ�X���`2p���LN]��-��R��d{JiΥ%�j�T�eS��[Kg��<�cI����gYE�ͱ�Gy	J�(���c�r������g�q�P6X�)�֎���W�e�o��2���'���
�h!�t{ʷ[�����ji)�|��D_p��2RZQ�ޖ����K�����1��s�Ʊ�_<Y0^;�B��rF�Ui<�.h9ʶvׁ�O �z[��H�ue�������@!Ʊ
��������t�����LT���U(,�b�l�uZ� Ӳ��'��S��D���e�Y�by=T�ʆ}M��7L�P���^�D�d7y�CK�7�-tL�s������*�p'������;�&�=�_p���%&g�z�]��HG�Ի�"��O=����E7<�쌉 R8�<�xWZ�;�S1��Y6;o�L/���^���+�4<�|O��ʟ����-��N� �(9ߖp�0S��vH����5�z�`e&������_j��E]��s�<���/�Ѽ���o�<9!I;���k�n�$��	~��J�5�os����'��Yz����O(p����J)�BN��+����iy��4�O��x��OcO�r�lU��'��3)��f��q,O+_z��������Df�{��ŋ���s����\�k����]&gr� ���u�8\y�I��۝�/�
���lw-31��c^���Y�l�kg��L�D5p}@*����'�C�>*�;��;���n���x$z�d�\��ރ�F����迟�p!�w���n3��N�jN�-��q;��--�X������
O@5�O�;�-�T����_�� '��?�ݳ�Z/Dd󪫫���������uV�Aa�S����[��k8�x�F_����B�}���
w��P$�ܾO�La�����KYpt_!v��`J�2V}���S`�Ì9�|�n�dkk����:wGf�ckѫr������r�>��+De�r���yr���ι���oPmz��g��Rl?������(F&8�Rן<y���]�L�P�?����)��%<�n|{>����.V#�u)3��������wc���*���0[w��H\��r�v�7�P⎟�u�x龳�qϣ��3���ll�f�F����������P3���n<<�{�>��j�৷�{��F���\q�o[�ך���0�xD�s_F���dV[�py��p�YeIx~��}L.{�c�+@�
��{�(-�]�������_�گ����U!8�=H�6�,*}��G�¤�5��72u�0��E@QY���%��d����C��Y�ɟ�VL��G����u
d�l�ɂz��FNm<���o�wv�Cf}��Q+��`J�L��I���c��
�����Uo�d/�=�i�4�?��m�;�	��$�ہ� J|�}�����5=�&Q��{�>$ܿ�K�����aݢ�~zN��rp؜i����hw��`��W	uz��&�dJ�^�	����9y0w}�,�ujj[��B�� `�U�@Co�����R?}�յޥ!lV��ى�����N@�̎+����f�N�T�k�k ��ԇ��1��^�R���
�z+�ى��Y��~Tbr�n�e�&x[`��j��!ڌ!+:2:Ҳ�>:َ�l6 �)��th^^���/�%�ZVɡ2P��[{��܌��q����FƝ�(B}�˪ߚ�D�����K6N�m�S�,m)<�Kφ޴�c��G�jl�P`����� Ս�zH�'�����\���:��%!7�^�A��5){	G�ͮ:g54�DI�F�i��䮍�,�s����5\�����>4] ��5^%S��̂9�k�\�/�~~��R\PbmTI4FA'm�`-t��3���˛��V�_��Y�_v��*��d?On��b
p�����f�ڙ,�yъߏ��u΋�0~ZIួ�_��"�W��ɧ�Ɇ��%�����p�&��p)�N�k�\T� ��L�Y�O�h�k�0����`����:��:����$���jݳ1�N�X��~���Ώ��q���S���hu��)�)j�hE(�XF\xc�g��d����I���TUB�o^�d֎��γ���&�4��tB�����q��=�4�D���q��;&�AfL���]a�&���׌�ǥ�����c�y��b��/������'�>Ѥ��kA��T.��a��m���mk�D��޲�#7���6d"�=Y�����I��|H��)�U?��\]���@T~�诞�2l��	>	�7Hє7�>��<
��R2�ܵ{�>���#4��~�`<��eq��+ O�U�����z.�����K�f^5�8�#���0U��}�Hř�h����l����X�M�9)�Qm��;�B@X�2�� �(���ut��O�n�X�SVey�I��x�X����'+�޸�1�%��'ՏBtXW\4��B��Y��B�ж��n߿
4m���1<`����{�0�l���:�Rl������=�b-�;[���� 16��Â�.��=���'�25--l����D:z��~ �t�+{�*�R"I�3t�L ���yo�n�"WA��Lrb��Mw%ŵqS�Yk"J8T	�����TH�uqTYzل4|�V��R�ʷ���N��������;�I۳�j ���<�P��Oؤ�6�	4ɏ �`�E2w�9�M�09&�5$�f� �/�x���AcU0=�KֿD7��Y$�T�,��31fZ�z�����G��T��Y�2����ۇ�y.֘;�/%��+���V?������z��cGPt�vɪ�f���E��^Jn�%���(��0��'�R�}#�x���4��+.�Z�i*N�7����̰�� }Ķ~@�t$j8�uu��s��ot��b����j(tP�
�����v���Y(CM%������l�A<���3���I*0����Ke��~|�Ě6;eXFHX�%=��:��0^��u��|�77���:�;�w2y����R~�}�=�J����/��9�Ǆ�&�:�����熁 U�m:3-99z<�z���,��I�}�3�d��Ϳ�l�D�_Α
��>�I��{|V'=�1�cEsI!�����SLv�=�Ӝ[<<ڎvksKdU�:8x�Ib� �t#I.���v���,���F����\�q#'?l�t�F���e�܋Jl��ȑ�`��JG#4�̴�w�����չ(�F��o�d�bɊ�2�PUˏ՞5K�а�N�� ���h�}����;�d�����
c����G*D����C�ڂ�ΚD����.J��:�(�7If��ZeЈ񽖞�`�G���z���݀$/T���k5Y�h�]S.�k��׺S�A��2��BS�����&Zd{|�@mf�p�t�c�7��Β�Za�2Y]|�kG���#��[�����k�Z�BY��G�=�Y�B$����?��rK~�@�g���]�9!:?���><y"I{��{��o*��l(������9����Z��[U5��m��v����)l5��������#�D[�/{guly����T�r�!Ŕ8Ɂedu$d�֥=Uq]���;���'�����(�c �?�
*��Ř��,����`c0���g�h{����6�J7�ZX�,�Y����Z�`j����/�O�J�B	ސn��NlO�����_�G~9vz�TQi޲1�9?���J��:J�c ��Z��Zk��@����=���;8Buz�s���yk�u�=�5�����2���S�5����ǩ�3;ĸ}�>t�b�J�Q�F���.F̊ X���°� (n����{*�M:�5��G=�������}� ��9����(iQ D��"�-;mu�Cgo�RhV�ߓ�(�9�ü�D?���vNn�̱$*)��k��y�n����ٓC���I����_uP��� |c��W���f1�/�~�@�Oy�W=�tg�J�5���)��Ϻ�=9��J�0�-���	��&ܤ!
�7?'�
^������O�.���X����R��1�ɝ�Ԙ�r�p\_��Dׁ�]ļz����}�S4N ��C��3�T����iL<��Kɟ�53��+G�����}��3�A�����n�2~͍_��ؒ�	��ۓU>e�������t2 ��Ƶ-�9YGM�VV�\e��
I�~e�>�2�g��������tKg�f�R��=��w9������^'��_ʌc&�����pL����<p�A򏧕2hF᡾ӳ?hg�=�����P��F�������|�:��<)JT��QT:�Qgu���ֈd�հ'�O����9N am� ;]�����y]��l��&i�t��px�t���a����
5E����OW��q9�H
<�k��5+h��>�{4�o/��Q�2rR���H-��2��!�;S�
~��f��d�7���ﲲ�j�n�g�
�~�V��+@k�A�駲uX<��gB���c��y�¸ǻ�y��C˴����Đ<0w.��Z8E[o{����[eC����	�<FX��"��3�?��H���_t��/����5 ��ޢ_[V��7N9m��z��Q@� ˬ����� ]�M�����vT���{�RmD�ZZ���hG�9�b0nyp��&I���x-�$�R��{��;��?����7@M�{ɟ�#�i��"g�2Z���5�f��\�d�\��1�pNR���7��'�s)�$�<�5}���ĸ6M��:Ĳ���Ѭ?K��>�$�o�IZ�\��E.B�jw�~�2�w�A�s^��z>T�8�s�.4�RH�S)�f�s��1Vso�`��]�����Zo��[ u����"�b�Ny�M��xΜt(�����P.���
/���T�&,��T�&&Q�O��(�};��fW���NR8�*��~�U��T5�h�p�$Q:۞&�3��c�݊�\A�<#�\��ҋ�}Sܯu5y�m�~�O���I���X�������m��]fΤRCw\[�I��br޵�z�Rr�����L^�*��׍@���iF���^��A����;��r��E�XO	����)S�+��D�,�����f��=R��A�`Y�u��ʊ�cIa���Y>����V.�XTt�Uu4�@m���)�Άh�*���$���t�a��[ź���I7b�|��am745�\!��0�!1*�f؇M� M�1Ԅ(�e.��"p������̢$�n��t�.)��Ϲ������OZ����� 9����SU--m�,��6�j�2�'�������E6{�<bWR��$TB����3c�!���mf�|^-ࣤ�{�yN�8���P��ռ\��ڛl�4�Ɲ�P��c��#�r����#��t�/�u�X5u�8���_0�9��x�tB�)���$��<My�tzbׁm��z��1\��o��y=�/�7͠Hr�������mr�2��c^x��˄.����ܪ[r�:�jYd��
�=�Kj/\��4�|���/5h��Y#���$�� �aZ	"�S�f����a�kT�����ȣ�W�ːj����&��� �נ�4�v�u�_�O
�q�7^ⱆ
�����ퟝ�j�մo�BCE]qmZb����_��0���t���R��-�n��P��Xz�VE�_3{�Bﰊ���/+�kn���-K;
|D_��X?V����6w]��2d+I�t��9��YG�t0y�U1)�W�Z�LcW�l�+�a*d&=�����$�%�������Ը�C�~�T-�+� j-]�L�e���G�/�9e�~��B{���1��3��,��?U���"��@Uq��>ˉ�����V!��~�#x�\��(bk�Y��W;R�xdU7��7�w�7�����CЈ�a���o�1)�܄̺�h֑4�Ƿ�"��)�v����2U�� q��^�~�Z���8tih��
{g��0�����яJ~�&R�3�&��Y�PZ]�/[+x��i��&i
�U�Z��:N�X2��.^����5���,�T7T����&�Oׂ�´lf:�I�f���N%�8�b�@�}�\ŗ3�]�ת������Y\Uf�1�b�k�A2IU����u��K��@�n�Hڱ��)Y㏎�M_��B��"����z�Y;���;�9J$#��%����7�W���V>5=a�@��뮉I��Q�ba?���[����z�x=��{��
p�R�X�p<�=-`W���+�f��k%�ը��8����`& 7�K|6/�a�u��u&���{h�Q�A�C��O)rV�9{���g�5	�]�B����<������z��I�Kܕg ����|�O4~U���Q��9�����*%5U����Q��JD�}�M�ζ~�E�0YB�2�0�Y�"����U3�_��0wD��.���H<��C�7n����r޼�����]����[���b#;��8~ Ϗ���G	ʧ���x^��l�Y�t
P��vZ0R�I��u0P�3�q�I��+P��Е鳓��;e4�R�|��7�)y�n��)Bmi+�b�p�����M��+��b�hS��(E?�W�@�2H�3�f��69d�x��T�m)quw��=rcW(8f��=	��saw�9��!v�ӕ�>���U#!�p��t��t�\�;�H�A���?� �Oյ�~с������ /:V ���!��	�� �M�� ��/:�K����er�	q�o��<��k����ʕ�m�1-�M�;�0��X��)����c�S�$��NO��c�V����,�8^���;TYc`���?I�l%)QJ86J�id��킧��%�'	/	��ǭ�t�˟9�L�p�F�B_�G��lx\��\�ЬC#��$���m'��vr��g�2�؏Lk�i8�a�3D�;;J���AH���p}�d���ܢ!tx����!F�Sv�/�q	I���8B�Q��K�����1��ܾ3����79HИ�[׿(�IQ�a_Ӡ�(��*��B3e��_	gg$a�@ө��4ŕa76nȏ-֙A(\_�2Fǂ�W��?><�ڎ%|-H���4e`�)���������E(��zw�ʿ �ϣ������t:�X~O�zl����|��K�	y� ��ǎj���}�f�Ȫ��9����Wt��xx�z�>�����>	�c�Й��P�4ZH�D��$S�Ӕ�v�L�+��T� �l�; CHe�26f������jH�(�=X�b��~i	I�A5�g}^*��~��i2�De+���Z�:#�g�Z�v| ��w�*���mm�>��]U��
F�D��ȩFG�c�r.���L�v�H�Y��Ҵ�n�$A˅qy"o�5o$k���K�B�m��<}l7��+.����O1�Y����\W���d�ڕH9N?m����]Ԣ��o��� � 6���E�¢��S����9$��=+Fɟ�G����;?���ݱ�OZ@�ˤ��5E�����B����]+v�r��;s���=�37��!\zj�q�!V��Z���� QAxw�{�fv��k�<h�C*hXh_����~��ס'�w�J��ì�Wd[�?�� 1=(�7�g[dϢ�6�p�j�|���ܵM�#��抭�f��e��JKt�,�j������ ㎉�R������PݐFu<(	%����҉��!!���`^��^+_b��/ժ!c���Q8�٭�Ns��P`����X����?��HR�+~��(�����s���ruU�`F�q���of�D訰�hJ�i��'iә� vzVA�돾�e�ȡ[i��n.Ls�GZ�_�u.�eQ�}H�Y������#����~�bͦ{B�!$v���u���<���m��kSe����{hv{����M6'4&F
��_�]�bg.}(AR�����2V�g�Ũ��ۨ���T����4yQ�=��yE~&�[OOl���'._����'輒U���G�k�bI�	����ֿ]�7�Q�F�D��8_�+~hS��>j�n__�_B�x*���X��{��|��
W�G+բ1��䕭$pQ>=,漨m
0���6_e%cbsP�t�ix��	���Z�c.dޢVk�p�t;�����(�#*��Bw�f��+I��8� "-���L?J�O%n1;���O.e�㭓E�}kr3�	Ð养Z�E�]۵�E��!��u�Yl���*/pvd�|�����Uҡà���*S<�Be�Xۓ�@�+�zz\��?�6W�(NB������|�f~Dgd�6��9�-�Ф֬���2�b�;��tĹEl��O,���NI�8ZLH@��w��f�H�4��j(f	(pY,����
��e��b�U���>5��?
�a���o�jYK8:ݕa?�l����l;q���z��G<
8�<�JH����,��!�z��&��nvV/rX��r�i�(�.n��N��RT�^N^J7Q� q�����X����y�c��v�,�T�^rN�F3�J��j!��9(��Kk�k����,,(�G����׫��	��.Z��D���(pPp�(yܛ����h��:5v�;%����\�[J�Y�z��͞��F��>���K�e�+b[z�U��L�������[ぞ[+�78�	Xg
%��p޷i8O��UX'���_
$�+����ιbpS�e@�-v�y�Hq�>���tK/ը�-M�Rl)_��w�D��G���3���� �*DC�dX�i�5�}
�ߑ��ӻv���@�������d"I���x��p,-e+�}�%7�%��t���@�M��3B:����/�2��&[�M�����ݥ�k��H��<��b`��?�3����4ڝ�S�6��/���[�w�2Sr��������i�������oƋ���l����~�M�S�Qɗ�.��$���n�*����M �c��ڳj�2��R*�)3�~�+������yQ�_�з���H`�	���C���_pS�znSƘ����ף Ni��~ee�)>��5�����Lp7~�\S݅ϑ��	�c==2�(4�  ��e!q�UK]����BX��C���#�2q�τ6�1��ץ�y������eFr'��eĔQ.#�d�LtR:�!�t��jj���֯�F�ʻ�����&T�v�K�-A��C�Ƽ@]��V�-u����`3�c�އ}W�J���C|�3e`2��Tw��T�O�����-�>��,򔌝Q�IT���.�[�Y�^�4�=��@$��ɼsk�EV%LɎ�4f4E#�/"�;�왻��T��,���L���>h�H��";�"ՓX�-B�d5��Bůl{�SR���^��h�� |\�?�u�Dȶ�L<Լ��
�%6#�h��he�*��0�VA�DMK�Rh��?1�I~�c�d��a+� ����3�C���m���5]ro�ی����F6�ہ�7��J*7��մ�A�y+��Kd�;�UV��:[���Cv����[-���l��6Y���q@kq�;.�ٿm~�C��V2�TL{&�(�5�i_�CH�Q�`�znx����o}}���'�� ����R������q���Ld������:��r�Q0��L�(�á�#Z�T8�Ax��Z�fߴ���
�d��]��� ����~.>]A����-��7əx�?��8^K�C�	�^d?����ٓ�1Ɵ�>On��2]Wa�t7�v��XC7�%����m�p�Y������K
��B+[S�Xhp^T��v==j	,G5��K���Ȼ�7���)K��� <����;i��R�f��׃`�׵����BipK5���J��"�UW�xee�
�K��L��J�m��'7^C.��V6�������rAzo՗���3W�[����kP�p�-� �/ϧ���|�uE�!M\7���x��8��y?C�G�����7�"W�֢(R�@[�����s�Tt��O�3�o-�v�.����?���c��W��ixz	�j������ŖD�0�V��n���R���<��G��O+�8�>��?J�F�a}ZV���b3Y�g�e�uA��������.��@��X�_0x�������8�tZu���L`;o�f[���_�Z������7�s��lf�m�s
��u�ض�"�"�DF؊���z�kK������dy��0E��(������3NE���F-\�����!��@�K�u�C�k5�%cL8I�w��W[��:}��֕�]�>_�����&��o5S�j��\ƞ��}���*L�X�,���&����W�FFg/�≛��+ywH�v��)����syĖ}����x(�1`��c���m&
�E��5�<�6xgL�����8�'�2�7��kC�C��:�R�u�_C0�{$=��Y�3��T�`�9P��ĀGd���h�'�a�D(3J�.g���q�^rn�}l:��Аʽ[���%Z�#%*�!�~Ҋd_��b�?xT�y�-|���N��J����+e����f�c�#�(�tP>:�_+u�~U� �ԫJ+z7���<r�:�1��v<���1m�.x���'�	z�{@�������)q�ʘq�B<��M��J�H1��O9�"�i�=���^�L`��9��������_�	F�>'?����L�W�KЯR��T�w�ק3�KL����=��ոI���q7D/�߻�~�Oi*p7L{jJ��0�pTU�OMk��`�p�_��������C��H��@V���rm�08s���!��WP��-%HR\A_����h#�6��Y�UR�����#�+e���C_����bu��@��c��[(K���GШ��M-,w��7���G��z�o�N���N��(x�:�}$@�,�%��B��
�V��0n��uBG�#h����\��݈�����zV�z�Ks-�<�QGEr���Y����_�b����(����{�Z	���G�@�263�22]�1�R������d�Q����732N8����yq����E�<Y��SY�B9]Q�6�ua�(�!d+�n��c�W���~jr&8�T�y\���E5o6��0��D��nd��4�5���'@�D���Jp �|[��C媟΢4�8��fYV�H�z� ����X�~�Y���!���G�mO��Sx�U:Da���3�s^���U�a��i�qq�Τ��r��jL�Ī�$܎hT�v�J�g�pJ��J�f�ػ���I�АL�oϻ.h�d�p�r�	��5�j�u�Q��1���E�&���\��N��$W�[�E+���g�n�`�W\؟.X���c�Z7=������^��M�uJd�Bb��{��G[R�9Uڌ�a�����g�����S[b9V�=�$��#Ѧ���CѸۋ�w����T����_��gD80 �_NNm���VH]��q��u�E�޿�#�D����q�P"F���P�[���
ݶ���L����)Ӝ���7�n�J�@��Ѕhb+��wǒ�����A�0/���#��?��:q!�q��u9��o��yH���Z*z���'[arڎޢ���UA�s���hiI,3���/Nr�&-���V!�oM�տeR�ra������fz]���~��B�QJL���Lph��=9�P*���T���އ �ߦ���&��u��Xb#�0u@XلQn=@��kCUV�9��S��y)[������G��iS�6�9��`�a�َF�ov�g�����X��Δht /�i����W|{���ѓ��U��O�`�t�Q�@<|F!j��ڶ>�@Ql����I��O6���yN�
��V,F����b7-�6�Urlڡ��Ș�bl=����2���)�0�)�f`���B�?��)��A��Y�bܯ�W���ܜ�����/�E]�׹�Wu�Tʓl�{yr�.x�����_S�d9�q�	@������!U�lo�rriZ�d���N\��o��j�A
��Ӷ�+y�}���f��.�𤕦6��P���4mA���J���8�o15׷ߘQ{����g��+B����f�-D���TuU��J(��~G�cͪZ��/�Ñ��*�w�

ȷӽ�3#{݇��El) �ԩ��P�I��6�U8�Y��]�Ԭ��u�7O#&F��Κn��x��T��a��Lپ�
j�r3-$1�e`�O3F*\��xk��|1s�j�P����)����W�9k�U��n��)^P!��;�w5w�{�8����ܔ_��=�t�pkm�?��ub�O��^�WSYv���׺�_��l�,Y�ȩ�pK%�U��@���-�PXQޤg��Kv��v&B��b"��Db����ֿ3����ן��X+v]���R��uo����������TQѤ�o�I�Y���O���"z���\��bF�I��DǏ��B�ژ����"-�}�|rj�����uX��]�Ol�o�ҁ&(���\wj19'��M�~�ൗ����{s��'qW���Z4b8|�<J�9<���X ��E0��3>�'D�t�If=���(_��D˵�>*���$�����+)X�Dɓ>N��goN����%�M�t����Ì�i�������`#��pYb��;���D�n!sdij;V�����_u����Ct��7��2��F䳦�4z��K������Є��gXTW�><�L,hb C�ĂR�EQDA@�h 齏�"
QF@� �m�H Aa�(�0 ��9�P�������z�"ל}vY�^���>� �n"���'�U@�ʾZ:v�%?��y��RP��O�WP��֎8`8<����5/�Η�㖜��'�_�a:ߕ��x4��"ںOf����{t�ݬ���o8�_=%�m��a���{�R)�ڑ�F���g�:T��(���b&������M��~]/��HO)? �-eB�C�W_���*������9t��S`���s23q=#�r��������E����M�:�W���d�<_�5��Dj�n[
�����X{&���c{�������%��,�oη�ǁ��Q�&�������;I���I�\H�w���|-@J�I�^�e~�Ț���F�5_}mi-6�'�o5Rג9��ۈ��Gm<�J�����d��x���,�Ǔ�!���ڗ{L7�ن��ʸ����?Z���&�����?���촡-_�<K�(_D��DSO�.��#,�:��]�'X�]����r%��ȣf���88�v��B����qX��PVN9��&������쩆I�0�}R���>���ށ���U˾E��X��E�5lv����������M%��eiE�ͫ�qgG�߁���cv��2�އ_5d�tD	l����ui���g�Ԝ�-E���j�W�*K���`�����.���S�/L[J�XK�d��o��� �6k���b��_��}5����� O��{��ek�d0�mW������=�'^�l��A��F��eo�5Aphg�Xm�0�'*�!]˞[�R�bd�>�Y�-̊z�l@��`�����}���>��,�_ԏ����gfLp�>�%�ī,�̙z�j,�ZA�/n�z 'Q�<��_c��eJl�hRIե���)�0_~x���|���=tl��ޗ�G��� ���]�7EZa��N����}�-y��:`��:[}K�} M�@�N�"��	�f~žڠ�;P���6}�}�4���/����ν�Ik�*n�+q�����=�l��� ']��_\=Gݽ%��/ᨹ8��F��kL�E1��d��:(.�w��%�l�M�� �����]Ăj��d1��fy��l�p�K��2.:�������U�����_�����w� p0o�֧��(Q� Ȧ	�����ꖼت���b��~����N$b8�nT��$�B`����y���h{�I��]��?�� �����A����3Պ�pG}�:�p���GŃ.Hm�8�� 4�F��+	w�VD������oF��׌!�.4H��3��{�|i/�S�j!V��)�I'�5P8fʔ�a�t���n�d����~.��b�X(��_۞����KY�)�P.��{�h4?�^���d��
�N���ehz%�pt?�|�'�EA�;Tc���M>��Y1���"�/�&&ZР�gao���ԋ�Hi��EL�?���DYc�;�f'4�
@ɋe�ɺ}�)�H������5�t�������������g���b���;�<� WՃ���noP<A@i�'��pbq"�jwN����"�[��ͳ�a��%���������]���/׌�����J8�p����K��F�����G9��v~^%�R���+�*;��W��N�f\��,�n�!ע* �_S8z�'��y���`=p(�b���mY����:q�*�/�����:�">}A��˷ѧ^�u��MU٧��4���?�M�iz�K<�~:��]�?E�l�,�HE�.�3�����2UZ�;�}z�X�����Gf7�K�jX����ʲk��	�3ypFx�|-������D\r[Oe���vԄC�L�u{�Ꮏ<:����^I���{(�O�m��9�yth�O>6�	j�~��Y��np�}�9p�0M|^��X.����X��	��?��(�����`4E턬���.�+O�{ ��V�VkBU�Nm��k���3��gW$h�ݶٍ�耤k#�� ��ϛE��޹����g�oVs�����065�0�9Xv#��O��	k�}��9 5W�Y�M�����.[��w���h�\r)�p]F��O�M^ �tw�A"���v�×�0#�P��D�n�m`M� Iz���T���0h�����Ur�HQp6��7�\wo�<�TB#�O��q��U6�����,��znE�_([�G�L�;����ǯ��N����paW]�G��	$ɜ"��%�;��g3~ʓ���K���eb{�p�숄��yW������(H��N�����p���D��ǧ�׽%��_���p�ǃ���|V�P�~��k6�/ݓ����?�ޖosd�5��'zڏSv�	]�s���v�����*�P��ۈw�P/����vן�_�zۉ%�`"Ur��h���x��J�݅I�K�vd��qw6	%�H��B�n���E��˚���;TE@�S�D��M{t<��I�&�V�����F��
����u�����#�J�����A�a
�	���6��N���c���k��k^�X��m#¹kǳ�XڂMBW��{_��_C>Q~/���K�g-K���� ��� �&�r	�G��������fzP)K��;D���A��a�9ɪH�q��|F����O��r��3�,a��3�"i<ǵdP�ZN���Hwp��(+_���=�����ˑ�7�oSqr���dm�+X�T�v����� �+�={5@"0?�+U��ܕ�,~�qy�
�,y����>�0�܂ů ��'�AcQ$]��ߢ>?)e��ζ���uo��,���kk@�� �Zܾ�����$R�B���/Yso��;��D�BN{������2Q4g�/������~Y<B��kO����GQ������ϧ�g߰:��?ڊN���q���ώ5��;��9�+m��yK������L�ܼ���n�r����R�D{������C'/�n�X�;����;����;����;����;����;��B�9�6�R+��л\���^���R�pE��͉K�..����쩝�L-|A�U�v�ԓ�z�E�b�'�%v��7���^�˭���{���{5�ސ�CGVZ��7l������]�#���gҶI$\{�LHw#ZY�c��YI�Q!���5x�H*��n�L����ZH������˓�2�F����H�݉yVf�n\���Cs��"+��u�_c31����1��59g��_К�o[ۚ�E��_K�NL9�ipTCz;6���s�؊U����չ�9�>7��\;�ҳ��h��Qd����T��엀�t*�0�X�Ŝ��>H��A��-g�t��-��5#��5U��ji��ġ}����ڶ��~700�Ԩ=ňgcx)����4�>�0�9����1g�,�,��Ф��ϭE�@eW��n�ų́�w�	��~^�۝�~�`O/�R��k���w�㛨ў:h�����ō���bK������:m�(�AJ��F���Z'�/���G|=N�̍���^&؍��/=7��Ԍ��^�D�@��r3�h�|��G��|�>��a/7�� \5������2�ǱnV,i�	[���p�# �m2�4�B��o!�����	��k��ԟs����;rK�ml����er�#2c%�R���̹�x����&*c�G���a�Ka(ֺ+1����u�-�D���^��v�z�ў�6[�٩��Z�}2�VIav��E�;̍�A���I��w�Qsʼ:��b��.�� �^ݵ�3e��p�թD��;i7n�X�pw�d�o$�NZ�9c�!+pv�>6
�Cvp韮�������y	�I�#��H&����VWt2_:��1����F��3�a$�Y�Q7�C��2��2!v�LW|� ��t��v�;ג���l6k�R`Ppg&d���φ[�:��������S;�xǟ���j��[v���¹�Bn�V�Z�l�dH�GG�9�82��ue�w*C�2O��p�3��qj;����qP�ZN�O3{zR����-��+�z���n�[�F_e�AO'��|.E��M�!n�K�M:Ag9S���F�?am�1�rN�α�8hNJ�_|�]bE��{�n$�������#}ֿ<�=�>�(�����ư�W� ��eN�Bz�F[�#���t{@�����,.sl�+Q�[5|#`���Vy�"�-���=���������ߧ"�=:5� ZX�$"���9�'�{۾���4J����nΗ?~�reB���pe#��0 8(�}��a��֩�وY����~��'�2ݹ�ΰ���7����C���|�餬f�抿0o��&�ٙk���[=��\� �u`7X����k���_�y'�>N�3�v�x�XH�I�����e����GK�ʿy@/uo�����pj�������'�_)7~ҋ��M*�՞{�-ӱ���������ý�䴁�T��G����(�z�c}����LR�@\�j��TK��LS���/p����������-�:~�w�����I�y�h�A�N,q6]�E�V�]����xt�ˀ��m"�/0]�T���70��5��&]��Y�
�|��&N�.9��Ck�mk�����dT�⦾Zց��Dh�E�ȵ�6�RZB*�+�?:W�vs�q�a<Un<�����0;�/q72��κS�Y��t{��}k!�V�/�k�w�St��$f��6�<> �pE�3�3���h�����Ў����3���Cu�[�����F��7�Gb�{ҀF1O�tmT2RʉM���Y�:�����]����뻯�A-X��?-l�w�[�ͻ"T�$D�+��.^���� ���T�����
����3�`�a\Xf9�=�k���و�^��@�*�Aѿ�	?l4D�_��/A��Al�{��!���ީ������n��Og粙�44B��	�@�3n4���jh�$y�������bi�:vƝZ/f�yw#��{��*?#���PAN�ӟd���KH�2�~5��ݯ��OJB�� C@+m��+�3S_��C�j�)��T���{��9T�=l�s��zK�P��Y�kՋ�����c^`�)��W�����b�]5Yr�C�:1%�6,�Ӗ~*���DC��
D�Y�Hj�o�_��xd���!ڿZW���	�G~s��'��a��I��NP9�'�h{�q:�h09ikg!�Vm@�=_��R���ݛE1�$y�&L�nu�3�=�og3.��A7������}v��kx�	��RL���E�I陏�i�0�X O�� Yr¯��1�¹�%��1�P��.|�}f�)����vZ�~�|�Z����ִ�*v;O�6h�vw�dP��5
���t%:�|ZC_�����80����Z<Y�A��e�zB?x�iwGX�7 B�yS�M�{ib�5�7X�@��}PS�K��U}?��
sd��4-���N������Uv��̼߂\h���A����I爙��N�)���ߓ��+0s>O^�M<��"��9���0�;W���#��фi��9���|�B��"���hL>�2`�E� ��S�A#�ؖ-��J������l�U{�#q
u���ǟ;e�x��A�l֠~9l{=�Um�Q��?a����e�]�͙�S�J��NF��D�O��z.�n(��:X���|�Y�M���>Y>�;f&��Xg�+�K"����O{d�ٱ_C����9�0G�m�H�����0ˮc�'m\K"��H���Z��f�/���j-u��ؠX���F:*o���3�
|J
�*�O5~�H��r
	�=�?Q�[���9$H�Bb�هC&��Tv��Ǳ���T���ֹO��c
�4s����/�fm9��з�F ��k"Ǣh�N��(4N�.�㏯�� ٻ�Dd�)��'�Q^�>^�ItJ}�P�;�^:d����.���m�ԯ��n�+Y�4 �#k�}[a�%Gl�Q�v�q�£�oY�REhc��=�q!r�C�|��[�`��Q�.����q�6Ŏ����o�q�-�O�q�)�3�H(r6���Ab<.�A�_&��z��˅���t���&�jBk�ܴҌ�?/_�v3�1���Wo�tѮh�<Y�zKt[��츽�F�3G�T~�_r��2�F�!)W��Ls�������!eR��c��n���p�:.Fa�S�=�/�K�F� T��#_ـ儼��w3�:)����3�j��L����)	}��"4�m1�:<9ܨ��ѓ)�N����Frz-4�F����J���X���E�}oh92{�N�1(����T\}|�6���K,αj��m����E��FUJ]�hP�A�t�k��{|�\�GP>c]�6���J�F�R��q�@n������c�}�{S�Y��pr���0#@ [Ef�][Ψ���G2ػM-L.�~�S1�u���]^�q���hx���p�nޮ[?�ڰ"�]Z���"\e�Yy;�f��<m�Zv+.uB6<���:6��+cl��Wy�xg�JYde��}�I���x#1���O������#����rb�We��.�=�/�<����U������m ��+�+�\M�@��o'���zųo��Z��19v)�P4��N,{�P~��X�r���c��e��ϫ����c�B^��2�p�I_/����©M��Έw7���ƙ�柜9�w�t�jA�L�o�O�3rm9�M1�-�\��NO&�j��X��oOx�L�o:���e0��U�J��� ��c�����}����{��QVME׮��Z����j~��k�\P7��FUM>�U=���6�H9Bp2kcu�*'����6��ߪ'���|!���av��v`�3��zˉE�P���5���i�Roْ=�	�&��A������#��ڜ_\��a� �j���cg��	%��x&n'ì�'&�O]`b��Sī�]�(
�(6N�c���?c�ާ#�9f�~��k<c�b���2~�b%�����a x���oS�bsŻ�:�!�z7Qǧe�{S]S�u�\a$4�Ӫ䔑fw��=cO�ZU����E����6|���
ob,��Jy�*{1-��}\�ݗ���B0Ҫ|�K��u���/��N�G&�;F���m�/uϫ��� �p���5�;�{8L�,���N�*T5ɢ��C��VE�j
?�������p��t��ޯ��_s3@�a0gR�79s��q0���v��V?��ԏ_@�$U�w����X8��3+����}������$o�V����AN������}Op���j)�g��B��������A]Ǽ�;������)��p�xu��H�~���/�H�:W��N({���(���ۛ��N��Cۻ�N��o}�e1�	D�"}6�(hv�ޯ� \����&�?ͫޜW�ܦxE��N����Y~HF��s�֯���;a�+7��\��Y :C��+rW������I'[�����i#��k�g�E`�QM��
q&:�
4�-a���\%a��i+t"����u�	i��J�h�$l�q�y;ӮwZ�?ڱXе���h�,�U*�� k������0?h�%U��I�|!Q��RT�����3	2��T��ɌšMá-�o\��+z`�'���b�Z��X�0�a�O�ݨ�<mzc��Gne�;c�dF����%��
�,�ыQc緙��5��ˎ����SS�bw�5_���R���7w�)1������,^j|�撡4�i��kۊ�9��1x\�o3O �n�i]Y���	��</��99��ƺ�gbL��(ur&0'�?��#;�9�k7�Qp �A<�x�\��=`R��>���beE]����[�2��)1�>r���.��_�W�ɕJ�| =����ޏG��j�f&d᚞�`���CC�T������8�#��t�V2��T�xv�wt�xX�q�KUE'8`��ܛj����!G�i���&?a���{��i},fm�N����F3(�و�]D�:�Zd�>��{Ã�;�	+rf�_nv7��F�*Z8��Z?S�@GI\��xȃ���`��R�&U��������6�8���O9�����5��%!W'���9 "�����t�	��|*���@W1�ZX�f���en\	W!�����Sl>N��s �t[�����M��T޻;��/a�\O��Z.OȞD<��9��0��U�<9�XR8;h���cI���E2�do	�h���D�� �n3us�ޓN�Q�F��)�I��U�"�����a#�Q5<��
L���I̡�����&a	��2��#���@����p��dt�b��w:Gz���8oº=H�M:ꉸ=�+� Q��!1�5�C��n��\O�0��#��v
��Q��+B���]���4JOy����==O�'U�e �\`b�[Mǻ�O'QK���3���P ^=1�JcxL�ĊQp�?Gd�m�wy��nl<��,1U���Hi���&��eW�m@��<e�l��X�j+38�[zSAB^@(�f�z<�]���L-��\y�{���C����M�����޶�gW�Y�$t��]�J�u��o�C5pvƵ3	����!��YeGu~��
�jά�C�*[�;��@��n��8��*L�fv6�(�st�7��{�R�?\���BܖԜ�f�ޛ�:�.��]Y��5��I�3gRZ~��t��������R�k	�j�8n\��E�نǜkl9�<�8hS����|Y�$%5/p~�X=-�d�M���OjT<  ;�;�Ie���	{�um^� K�x��/2�ᕹ�Xc��ԣ�rbc�q�`�ź�K�*O�M��EI׌�%ݻ����C�bT�	���B�vQEHr�Z�(��J��W�Ai����JE�%r���Y�Q?���!�&�UX#�1 �GWd�ťJ�߫P�����<���v��s�\H�vr�N��Tz$�j�&�7���_l�jdÕz��$& ����ح��q���N�o4U�s�qa�Dx�J<v ������@qo��d��NpN*�}�@��ݨ��s� � �!�D<��f�3L&�0/�U��f+Ф2��*�Վ�P����P�������%)S��ݳ2�N��*��XdJӃ��4Ω��z|�%ȯ.�y�΄[�,�#FJ����v)ԗq��M��*���K���B�?r�b��aE�:��ϼ�4-�Ï��l��6��U�A�.*��4�;tŕ�k\��feKd	��?�R����u���w��L	솨��I�������*��:�� �0M��ÿ/hN�����P��D�B���1՝��x/ɪ~뎃�K�%��8Z�u�X1�&�4�D
�X�Ĺ�S��E�04ST�đi
���� �u!��IS���=)rB���2$p[�758�[�mT��1P�����fQ7�O�C����z0����;�ô��?�H����Z�cĽ �j!�(��8��jTUX3��qj�/mHID��Ӿ�?Y� 8K1��0��d�;� ��a�������;����{�^Y�܆�K����Iԓ;F0�w\mFRj��M����������{�Ԍت!�������
{!/<��,���Ow�}ε�����-�9�5�C�
�>�LK����:��퟼��'U�`y�n�HJu�9�l�nX���zѻ�[qOR��2{ȓhIz�hb�O{�#�{�*{�H��ڍ�l��i���F �S����QHX���l4��D�"b;��3���ح�>-�f��{p��ղ�Qgs#��	ĺّ@�|��[��s���P�h���ȡ8�����P<'Qmv@�+��2O�I�wJ�ЇK� }n�����Ӌb�Dj_ݰ|��x@)�^���j�h]���%$��?�L� �7@�g�����l��;������sM�$&�D������������.�<�N�b�K9�D@d��0��Q�Вs�Q0�Ks����t��t��HمF�
P���Cn=_Hf7������=��@u��)̻	��T�E����:�kR��{���{C�#��H����J�:1��f�������T��b�Ԝ:E� eD0��~�U�4�.v����_����x\0x��HA�x���g���Lħ�b�H���Hl�B�������{x`M�Ԣ]E�Q�X��&T�>X 	�?׵d�+��O�b��5Z`�.=�mW4i�Sh��%y/�_UZ�~4)?�~����")��c���1�`|CD%oS]S��W���n8Í+i����N����-��J�����k4VP��M�H���E��`�z#6l�],�ݔ�ک_�����Ǹ��7����f3 �.+qvY,�ǵ��
�b���Ķ���K���P���b'��j2�@-ľV��-���AF�:l�U#b���+O���z�j=r\5�a�c�|U���kP�ͧ9�O1!B�.RHw��Y�T���r��.($Vp�t`R�wp�l�'"��6�\r��]�/�4e��3�$;NW��8�k��E�hH��嫆,�*��X���bJ�)T���7�������3C�Č;>դ�a�#>-�~����/�������L�@r�LS�Ѥ3Z���-!E|�Wz]�g^��A�ɭ�k�ѓr|1XG��@����rE��L4���n�bQ�;�Da8�H�Dq`d�,?t#D�2�q���Gy˅��P�B"SU#��ъ-��B�
�'b�vK<����A�~'�Y�x���bLM�"�p���4�/0�����*]�^��M��:��WI��Y�����9�|�7n���v����PlZ�	�E�)�����J�خh�!�.����u��@�Ƨ.BU!�&߃�g�=�؀#�����h��뎪��>���*�L����*g#��w�[~G�!�q _�O�{���y��!�#���(��]t��0�Jޱ8����Dy4�� 9�u v�W�$����/�&�w��k���,���"Ƞ��P'~<��	�9X��H�}ha��yɱX��73:�����x=b� �mF�?�y}��F�
@-��#�_IoC������l��`c�����GAZ���[�J�69<�ħ�����	bM/����=�&�pT��(�ina��=L3ڌtU��nr���XЄ8`�[TCSD�x�i��C���zİR� �*��s�l?��EzH`��4v!�=^����|�-�(8��oi�[�>q9�13��ճ�*ԙ��fe�3���!�� ml�&�ˍ��V�Ux+%%�8r@r	�K.�/���v0D;c?Ym�?��b�O��]�-�)��P�T����=��u%��h<���\k���㊍N�̃n�<��M�r��O�:&s;}�g'�_�ܧ��*�2�
�7���'�!�A��m�/fԫ���$e9���X���}1w%�I���1�О���Ze1�ʉw5��?�\D�,��!���.V���W�x��'���m�=���8��ꨶpi$ztQy�2�b�u�j���	�������n H@���Ć�T����?�A&ʙ������YC���Ƌ��W�[�7Χ��Id�i��H��'����
�Jv�_�+�:_т��s�N�W߄���2���箻?ps;�f��˞�_?�iX�{]���
V_�> ���"�]1RBX��|+��h_���Q좦#�eT���#3�����Wa���{�K��
��Ox�����9M�R�@R�.ު$9�L��ؘ���8��1���RO��1�e{b�`T���DM������-�>B):v������.	��T�~��t����.bR����g:h_���M1����J^����oa=;���7e��U�	�A;I���l����������9�x���mΝOgC�h����/�@��i�t�]T'�3�Yp)�E�ʳ���T��=W��0[ݱ��g߸��W�u6��5�Q�xSG�����W~���s����ݎ��ݼ^[�D����e�L���6�مOo�wk\���հ �H�8PE:M%g���^�V�~��n;�ݬL�*C��n�TNb�wL�~]�ޘ��g.�?�E�D��l��XRD?3E���B+�(3���t�w��y�a�
�[����U�x�g�;����sg-d�����B��W[�
~+^���b��}�I�DYH�p����T�,��f���=�+^̈��ln+�rg���s��S���f�u7�&��PnqX%��\�H�_�	�j�[�u*��i��e����*i,���P�O�7��(r�a����AO���)9�&�'N8t�e�}%z.���HUU#����O���8M���7{�q�.d���?~Ζ�r��ju�wy�E�<�t{��Ā�h���9#�I���]��G�;M2J[����S����)�M������+	e6ӹ7�6�i���T����In���	cnߌ�g����z<K���
v{�y�2��5��~t��!�hF,t��vN���xk���}�� ����A4r��n�ޤ�ӗ�~|o?�w*�H�q=���&�hh&��Pf� f>eD_O#����Ԉ��}����ĉ��w�!������ښ��3Sّz�p�a�q�b�j&~5������-����ə��S��h��%��w��0�����0�
��������I	hD?����,玳�N�-�1>�����S�Nhq��ʏ<�-��77|�9"�AvIi[�Ą��6����"|W��z\ko���W�ig��p`�gN�Ee�JͰnL����[%�I��c���݀��2�v�����^RzN/`C�qF}tq���	1bV�]�ճ�2x�2�<��)8Uʢ��ȼ�l�IXe7��D���Y�b��8��;�V����kR���ӑM��|t��� ��ǹ'�<ث�����5zt�K�E��������;_R�-0�;�iD؉ن�Bu1��8��tiLb12D3�bR��q�dh��Z�-��w����ƺ�:���^1D��eK�J��4�j�i��qـ�B.�����A��Н\+�XJ��}tH����&�ﴜ��D�JM�4�Q�#�A�!�Ik_�������Z�ҟX�k��5#(~��V.�=q6��D�X�aR��7�l<.<s���jeg֗j�H]�a��a��S#e�m�����Giq�{��4�gΛ�|��ȧ�8�5�]6�O�H�aN��ե�F�iF����){<�o����'Z\���8<%��L%ݓ�'��G�)J�(ă�NSN���s�kxs����M��2�_�RǦ>O�̊�3G�JC�5^_������7~^��S|�A�����hj|8kب��N_��i�3x�>^�ӕ�<��W�y�2�a��cՀ>�~;u�ߎ�B11��85w�1%�k���z��-.����q��x�@.�7c�}��P�0�����\t�_J,���g������Φ���~���ZCӭ��3�[�$�f$��ˆm��S�2��
	G��g�he�uk�?�.oz�<e��V��Y�f�}�l����Q�r����Z�9�t�ԥC���:5j~/��Li��7��X14���N�U���8K�l�����a�D��^޶�ja�z����Ϩq�Z'�Q������x�0���,^�{��>W1.O�s�3a�;$z.�L{sB[�O�]����Jn_c��D��F��N�c���dn;�s��i �$�]�D��t�3?IMm�5����'�V���:�C�b��u��޳O:��f6��Zd��C��E�*UD����\e���/ic_��#��������W�w�::n�S86����U=�[�`��M����'nz=��;������Ѭɜ�U[Vt�;+�h8*�W���6C/�O�Y�ki��y�)5z��H:7zK@��~����sgL���)YO�<ҽ�
X�7m3҇x�t5b���g�H�r����x��'&AP��ӎ<����TƁ��%�[��v"xؕSy�uiI=%��/�IQ׭���7U��,]�v�_[&�N[�j����F�&�;��]&���}��T�͋�g�r%�^����mf5g���҅�6������p��(�������2z��_Y�45s�7�iތ7)����`)fܙUV�|v��=j�it��v\�C͏oj}_��v��.���Ok�{L�59k3ئ�ڣof&�x�g��y?�Ꜥ�^��qj��.ѣk%����]u�<�ˣ�݌wО�i��%r���܀���	]<�n��GT�~'�'C�}��௉�Y�NcA��p3���l�^�?�G��Tk��Ӗ����i}u�W_��}ȇ{�K/fS[�^Td�����.��gƤq�i)����6���O�ǔ�jA�v����x`��
�F����w��4�׫�L�Au��Z_�TI�[&��{r;����C
B����i�dٴ����CXu��)f!.;vX�n���u�W�a���T
%�A��0B�mmu��A�|R*L�+�흖g7B�QӔ�'v5	&V$�����ĸ���P|Jې��N�9���47ϭ��B�"82i�:z��q�Ln=1��9>pI�ً��A�ͰS1z������#���Ǜ8�P��>x�X�t��t�Ha�Lh� )���#S\ǈ��2�����^Q"�˞��1߷�޼�����	��}�.�Yn���%�^��d��FI9ھZf�ս?�oݟ��1%�(jk����w�sN��Z~�����HuM�!���X;}BB�Ւw�?LBѹ�xV"q���7�.R_&m]�	�z ��J�HC��f��g_�cB�=}�fH,�Y�;nS���`1Z����
��i��Qk�m������`�X|��c)�8RtM��M�D7����qW�6�ԫ��;����d�ѺO��cv�v*�!X�}�����>m���c|���zeǌ����C�Fx`�@��� �3��Rқ�L���O�T 7�e��@�H���j��,%��O���wN�􄑆�[J��ќ��8_�a�vwS[��r�� P�w��O�n$�G�|P90t8:�y�����׽ 8迪�Ć��!���;?��b�
i)���d�Z_����1�r�T�i�pvӴ���/?�@s�[�'󴴟f@Y��4�G���hJC�N� 8��Qn��jd~����0��gM���!�H�6�ޛ�]w�y��7'�#Q�J㾗~�U+cf�|5`�Dt��nN���0�� ��j������@h	܉>�2��{�ĝO���c�-���k�Pa���� 5w��B���9����ѓxG"����a�~�l����X5�Zp���>�$���'�b�w� �~�5��w�^�72N���r��,�L{g�� �Z��z�%�N;Ih+��M,��5��ZE27�B��͕I�hH/"��9���t}��b��РbJ�y�'�A�ɣ\эJ"em$�'��!+Ox�D�+�x#���m�zQ⸷���i�Lþ���<��~�0��U����P�*q�+M�o���*gAOM<mکA�Fm
�m
GZQ����}���#��=1u/B�x:�L���?��)I��CYA�Z��:�쾮����9.�Ȅ��x��U�iڊ�R	�|�$��:� ���O�6]xo�߸�Ï�|F�SYF}��w&�Į�7�N����XW?�&����-���w�}|�9!:5tLc�˭�4�3:�DY�X�OSs���d�z8�(����@�~Y��HiL2D�j΢%��b��΋�I[$<Ɠ����r f�o���M$����bD���Py�����C�r�x
���ף�� O�~/mJ���E�'����@;����-��jmN�į�B(aH���V�2ӵ�Z �:�a48���c+n���!�d�n���WD�_�E>�-K���S�-�:Ϛ��-�����	��(1��y�S����bP[sZ�}"�Cщ"��wL ��w(�`�0��o�~q�L1~e�z�����i�𴓎"��(n^��%�S'��_�<A����\�Ͻy��?Ag�ヱD�A9�^S�G�:Ju����RPұ=غ/�/L�s�����L��4�CM��� E��ɧ��������K�o���PDhHޠ�'��|��Rb�}�{,8�~s�wG~��g��Vd� �nRp".j�麙�ŷm�L��ks���������o�)_�t�f4Ppx��O�D�=]�f���K�H�1;�b
�y�|@b*����r�Y�w��\��������!)�Qu�PU��Cż��:�K���:k�?a᠂�
Q������m��[�^������oy%^��ﾚ�Šzg�h�_'�����b�-� �y9��,��o�[�͖H����l�·#-A�ߦ7i��9H� KE�hj|��?/�?H�]���x ����{��i�Sa̋��_!����J�R�߄��3�(�/�%�
dI�f��/1h�3���
'�^�b��1���L=��S�C�Z��L�-@]�F�o��݀S��8EmJ��r�nҳ����lZ��B���1y�cXM���A��qn�D6
O�CK���䥶A�]t�;������߇*m�"�lz���ܥ�/)��׋�r
DU�� _|{��?j�7P��+7Cf􀄅�HT�]����4��~�qM�|R���2
�����P�� �-�zu�3�a��х;�y���-z�M����QP}��Eڀ'�������$;G�d�_�X��A�߰V�f���U�Η������2�.P:
*�;�%��I�˨٥i��bZ��X�Vޠz_�r�K��6��1ZY,}�#�H����c��]w�3����	R���/5s���?�Ca���6�b���%^9~^.Jغ���-��K��1*C��r�'��?��d�|O�����G�K)�F�'t�S��ρ#-�ߜ�!{���9��ȇ��(n�)WE9�6d Q��"!�w���ŏ��!�Rɞ�~u��qv�¿�Wr~�^�?n��X�4����Mƙ0�D��Ma��죋���p&5w�Z>^X����.�

P�����Re�j,�;ӘX��`�1\M�l�p�ͥ1ʙ�q��czm��T,]���$z�F�tN�>�η����R�]_���/�1��fw�\xUzTN󕓩4�=��Si�2�>�L�E��  �$j�Z\\d�kpL�S)��5�G��&q��%*Ei*H�<xme��+���vI]����Ћ
��n�D!,���|���X�XX3�vo@s-�׉����s�7������C�D@�H�
[?�G�giP�Y�yq���Przs�������M��:N��2�`�b%p�_�`�1����P����^�.�uH?�����_͍n����Qvs�m����HeJm�<Ԓ���W��y&��*���XH5��x*s�:�v ��u/�� ���BA�f�ț��H>&���"�\�[��6C�4�_:�8�mn���"C�8�V�C鞎�AG����E�dSp�sl$j"�X7p����X�!�u�W4j0���SƋ�C�t�j/pHã/���'P���?~gR/���#(�τKǻY&{���9�C�(7��_W��-NB]f.�X���O�4�ƧF�,�	�#C�	�>���Ρ%5�6ɋ���.�_r��K�6W�6�8*�ӏ�[��c�&��UK�'��y�]H,�� zb��;��b�a}[�ԜG-p�z]��~fڜa7e;�C{q&���s=7�-7�]��ҷ�g\�
ϗ��hR |�0����#��6�A:�Љ��#f��YɊGޝi���>.YB*h�g&�vX���D�
7�3��+�q��)����y'$)�4�{�E����`L�Ʒ���26;����R[��� ��Y��C�ݣ����RB@��v-p��:{*�4���_����ct�K�-q;��Kw�UA�D���ʎ4}�?�� [9)(j�JI�	 !`�.��i4���MJ~
�/-�����e����;`�f}�@|�Jm/{� �]��Y�H?��7��q�  H���־���7�H�R�Q#��.�ɲ���2G�=�z�ͦԽ:�/�@?��\B�~�j[W�Tж�$�3dnKpϦ�RNH2��¥~�TS�q6�>9}g��;9c��浲{u��3�c��l��)�P�s�~>7�J�͜�-O�z����{���\.�&�kw2y�����/��*8�?��>���G��?l���t��G���6�D���N��~H�����<���oKCy�5�9ͶMu9j#&H��6�FU���Q;\���(^�>+�-������i?�B+Ruͧ�I���X�n/�e���\�k9U.�yin{]3��d����D<opl5<-<��/$K���'y
��-��_@|��vU+��-�<,t�v����{��454TO��+��։#�Ɯ ��'���5�C;����(�*�v
	U��_p�/^F�Թqk$��
e����q����/3 eD�9���f���d:vZ��m���;R���}�]^�9դ�^Ȥ�5Ri�r?{�#�jؘgj��X�ˁpT3{5��|z�H��qenZS/�9���$ˁz6M�pL��ܸ���nB�\����N5,q����V�][q�vu%8;{���%d����bi�����^�J����ڋ��~(4Խ�x)�2�J�quLm��v�)Ԉ��`��^>��
�w�;��m�d�t-8S&�~�n�Ƀ5��E�>"? �?���%je�Ԗ��:'�$dHW��Q�N��>�:�O���C_�xb8Y�n,�q/m_Jb4��>1����R��W�n�ժ�N�4���[�p��<_.|���_I1N�zҨ�����-�UW#���Dee;����\�s��`m�B�������yt��qm����6�
YөaW�N8⹌�nj<|�ʧ�M��T�.z���Aw�n٩S��Q����V�G�V0�n��»�����d���T�i{"�;��ߺ�t��b�͌#�i�Ƴ�ۺ̞�H�� Vn洞��R�K&����ǃ���MU
+ٛ�D܃�o� �K"�)�c��4e�<%��p�UUd�Z8b�:�1�%���<c�[#��������G���<c���ItB���E�*�u�����+'\ E��磞�V1���.q0����=x�ў�����og5�yױe����[�:�iI�9�$��)���(�ˍ��~�v�9dB*j��v\S��C�⪇+ﺪj��ƕmn,�$#G�y�� � 4.�m����0�sa�2RvPU�X�k����<�����:G?�p�����<=��<�k�<�87�������ҫ1�@Ч+���v{��ԧJ&�{�y-���[�[�׻^;��%�X��~�s���U������\k(^���O�+)Ó�����J	6�0�EՃ�I]/��o��z�	�4�v��u��~�#Ovq��?�y���j|�S%M�;Ŷ��9uD����1]BjjaV�sB��(y�!G����x�0{��j#�� {�m�O��nt*���B�˼S�5������p���L�WӦ	��"�r6��"4x�����������J=���)��T���Z(2aZP�ٙ�J�Ǟ�bHJY�T�^dO�=��;�w������>��|�����?�Ϲ3w�E����s~��$H?t���b����3p͠[�C|�R�n&����ϗrf����#����֤�Y�'k>�t[	E�i�;k����{o���z̶���LG�zx��3�`3mQP�g���(kFڟPQ��{�=l����E����uLav�����w��=E|�\���0>�V��]��� t�>�i|RQilŸu^��M��� 3��5���H����W�Z$]���#�{:����a�_��.�S�[��'�L��� � �ׅ���t��^7/�P6f��Q����|�Z�	�/-/zn�N�y6�a!���`�%���}N�
��]x0�ňP	���M˛���~����ԭ�bD��|�����/"�#>�[S��7�I7��v��l����l�^�d�?`���J��E��S�Лα#f��y{ 8(��	�_�,�]�B�F�۶B��c��+�ߌ�?����<h���z��
�u��}~�&�nI^���L�٣U���ߚ�����s��RS�I]���{'ނ�K���җ�i�+�A����z��Y�:��C�����	%��w�K��kv����h�0��	T0�K�\ҳ	 ]R���)���ۈ��P82���#\o��Ex�m��2��z��9SajT��_I��m�B��js{��б�[�?�����C@y>?hzlb��g�U8y=]�T�~��<��	���u��B$���\�J��,�gb-�y��0'o�j���O�$�Љ��~�u� X������'՘���|����'�г�b+�XhD�)�ʯ|QZ`�Y�� K딓�6S`���LJ�z4��Lw�8�i�XRC�yQ�Ά�l����K?���c+;#�$��y��A �b��P��0%%����������AI����ATsQR�&A���K�[���
 ��S�EW����l�ተ���:�Az����aM�b�����^Iv�У�t"��&}��X1��o\�Dd׽A~P������QK�xE��G q9�6!�+��V<~����&%�#��S��<�0���a��6�]i �`2��2P.��Y��j{�I%F���Byվ���]���͔8 H��lR@ki�y�y�!󋜚C-��V��t���>�e|VR�yh˹R�x���w#"���<��<�����v��7�$hӍTr>y�_R�t�?hn�iܫ
,�F��5�q�4�V�l�Ƣ.�U&+��Y-AZ�7��F:���6�_��c^1��u*J�x�z���V�<M��
�������!�S����Ψ���/!`\u.,9��`�h_����_�";�K�}D�|��E~XNe�ê&�������T�������a�N�-�P��v_R\N��ܟ���e���
R�r�DHG`&�oJ6u;tTt�=�&��+�Η�@��}μ �g|wV�3��5��x�����*P��¼���2�%)3VC_������+ѹ�AMKa���s���2t��7Yee-��f�և_�bL'~�SB���ڒW~�*�[�`i9�qL����ҍu�b@�;g�j���#��쮈1;(���-lc�8)������\�N�aj0�OJjKYH�\�B_UXL�Á��ϧw��r���N���r�=�(("�u��k(Dm��b�K��N�@m'*m]EY��TUk�\�?^ԕb�?��X�{�R���+�FX�K�Sk 3q]�?D���`��T.l'@Y�dc�q����<4���m]�=]�+�Ʋ��FV	+��\lx��3������l��$~��4�I��@�l����b^N~Ԇ��1,�z�W���1Y�hl�j�Y����E�:�V���y��?��	���-F�y�A�4�<޺3�ﳟ��W	�^5^��;��`�l`�Y�	���?������y��ZE�9c�)-<�f~�c\8]���$|SE$�\�>k��#���PU3����Q�n����������A�S��BcQVh��I~�3^�4��5b|Z�~ �\c! <�e���p���R�������C�O�~�9IM�0_*+��u\���������"�YյH�!u5Ξ6E�|�Fb����"Ҙ��{���%Q7��ձa��VBmL�ɔ��MCT�0U���:�2|m��' ��%1c� ˵+>/���ޛ�eU�1���vv�T8��A^��P:#`���N ^�R�*�$� ��?ő�]���/ރ«��g:�[�u���sm>8 6 �Vt�"��>|
\��&����l���m���� ���U�ٷ��Yl��2��P��J�٥�nE�*��ف���	xRb&�.�@З�/�
qs�cR��H�f��������V��F[f�.m��'�C�1�m}syq����d�*X�y}�n�=v(����ї�	*�+Ũo�,�G���
�U��Q|D>�_�{Q�x�1V�#�Gٰ[R[��]!�����<�o�y���&�y��K��o!tN�=3�W�,�]��G�������|�*�����,]�equ�����WvhK2�8��U������ma���9Kګ��g�m��̍����DWn�J��f���0)��\�S�mR�u�b٢���v��L.�,}�X�`��_T\;�:�`�X���%M@T�Z<^U���5�&~�\���@�F�*{��nK%Fv��7���1EڻO�KP��7QA������4�ڬ��u��>׌�L�BM;c�5��|Y��Ľ���S�F|!�"g���@ꥩP5��3�vn������ro�g��,L�,9�DD��l���>�}�i"��Ce��N���٪�}��VPJ3�A<ѭY���ߩ]�	�����F��l�oG��w�i4���x�*��`�!I�V2��Ï��i&�5�|�g1�t�5]��3v\=�#�c�����@��ύ�E��hV��sޭ̸�g�nWqWūY"3)m�qm}���*�0k[��lB���1��=]i�*)���|)�Fti���Y�����{s����H:�ژ���l���/�3�L�����ըx"�
�?c��V������_��psd�uy$%�׫�W!���)Lm��C�s$%ň��}�q��<z��y�^��(L1zl�r�ӕ�� ���ۏ=%U@�9����m�הּo:��$�Ի�����W��uд�����a�`Dy���,|��8����M��*��cIW�0��.D
��r��"��Ct]n�<ba��cq���8�1m�yܭ7�L<�C��2�d���(�@�ׅ]�In��f7r���V�+v<\�$H'��0�י�[|�_�/�z��78�#���=^�T��ű�aˈ�r���Oa
-\�1��S�=�7Mu�N]$t��M��n�K�]E���̂����C V�o-t-wFg��\ي���I&�c�m���=fl��A�|;���/��ʰx�̈́�+�G(zDZ����Ʈ�!��Kym���G�7��%�"J��lw�����^�,Z(�ME�	���c/]J��I�DX��:p6�p"^}�[��U����a?�����u�[*��.�+��L�/6��ի@q_C���N�`����=J�7�_r�j��j��̎�c�:�������Jj���N���"n���;�����v.F�K���FW|<��K�W���H�}��:���� V�����&����HXGRd��-���m�0_���HXF�)�f�M����kI1�J]��;�w���u��T,ў��n Ԓa*��! ��7��:Y�ԧ>s�-�u Z�+��n�*>nn����v��	 d�%��K�h��ߦ.�l�t��#g�I%���*C�э�f˖��4�y�6��iE�ϡ��w�^	cB��C�V��O�ˋEm�9��� �7��t�>����9�u�����A�Ins}g��������`�С�R�8�&p�҈p��qхhw[?t��io$-�I ��W�JxlB:~�>��oj��~��6� 2T����O}��++�6�����m籟21��U?�Բj a�^ځP�\"�Ah���&�_��*��u�\��f���=�79��b�W�T��֠�S\���_��]h_������b !��8��j�@�Yӷwƺ.qx���;@h�G�Z(X�NcTI�l{\2�@�4t1?��y}��y��@�Dn������N�I[�7�i���h�z���/GPO�cߜÉj��HSI1���,�^�
�ng�E[Q/�ڴ��ϻ]�[����'�Ae!�{������nQ����w��iIc��F6�gj�H%��Hsݐ��ב���> �2 ���!�:�FR�Z��2?����C�Ŗ��� �>�K�G"�G�$�;�����hg��lz�]�d�b�]�6a����c��KK㖋�Αˇ�E�j�[�c�!��߄����Z��ŲZ���FƳ���H�OױE�#F����b����}�_9G;Ń󇾚�Q��ߚ@�IY��mU �2����yhK+�!0�mv*c���e�����A�?���!����Nי-�_2���cCҀ�{w�����+�ed��FI_�B2}ض8�{Bj�)��.OVIB�=W�gO�5�A�L���o�vL��/D��n�c��t2��^Vk�E=I�n��nש(6um�h�/z���>B	2"�@�,Tpr�\c�#��ʰW���$zt*��Qנ�lfatO��7��&���G��gl��|���M����pb�h�Q N2-M^B[��T<��KP���B_?����y,�t@��s����+��	��P�<���j^0��#Bv���_!���ā˂��K�Ϡ{�a�M�Y!g��=�L�ʼ�3_����& �m�}#�6��,&@2��*˘?�����-��2b�Q�HghI � @^V�j���D@���ר�)���_�Z]mD p������ ��sϰ4��µ�����+�s��h�/pr�)zч��1RXɎ�p��KV��^+�"�;���ا0�ǆ�n�p� H��c]r1���i~�T6{�Ģ����☖u�j+#��[H�aç�OH��譢x�\d���Ø�|^����<M����u���s��r�}��~�[ƾ`�E�Cf������k3v�*�z�t�5������J|�#w��b��W�4���>�g�3���w6b���}P�Of�������mOqX]a�^�o	4�`�⤹/J#&���@F��:	Ҧ��Hv]{ꂲ�M�����0�s0�?�ȓ�nX�ex�>�E�j��Ȳ���ai��=���t��/�Q�A.~PY ��i��3�FK����j�a?��r6G�FE�lފ1�����'��n��>�Z�e�LVB��������Fg1\weɶ��RY�6�L=�6��ʖ�D<F��Ff=�  T��Ā�#�@����/z�z���T͏���^�V!g	��̋��d��~�"1�np�x�q2hH���ԩ�_��i�$F*��όD|NWx�<�Ѯ�(�L⃘��F��񣚄��64����r懗�W�
�:	����- ��<2�i��14��[��� ��~^�Mo ���@��O���1�_�|SaO���Q�����n�*HRؤHS��ѕ� �G�[(��]u�E?�컼���:�?z8����.H���הF�ɕ?ڷ%Z�]���d�`�N\&�`�&��ғD�Z�FP��ʵz�����W�t��!/یZJh˯��+cL	�+{-�]9Ni�������!�v�./��
D��T�����a��@h&�ۦ�`j`I��z���%�7f�&z�k�b)���}��| L�H��ň��-�Jl��x�LIf̧��'z*Ǐ�.z�����?1�C�o��>�5�3�4�E|Dq��{�Y�C*��d^����*�F��d�		�%#���\��J�Eñ	G�?R�g=]����%�����ư�L&���!1����spf̷��|�^�m���C���c�^2[F�VF"%{�9#��)'��9#��h���/���PE�vn@��t����_4+�W�sd�)���M���G�	-4�Z��í�;{��l8�щ΀������~ʄcZ�݃\f��c�ܠ�]� �lBtY�^�1���C{�{�2�3�.��j���jYۊ�+=��!�/A;GS*��*��Cdf��he27��yx���2�Z�6���k�G�g�Г��x��Ht:}+u��ؤ�/3��49+�Q��V�ѥ	�� tR1�0?{BF�|~��̮�w/-}_F:�6�����Fڏ�R�=�pD�7�����n��=&X�r��G���B.F�`Y}r��K�v0oy��fgg�FR�;?O��Z,���Z4����e��6��q'��-M�7,�H�?�+�
H����{1Y}�z�o(5�׉��~�XB�Z�j���y��x��2Ԁ��P>Kq]��_ rG���t��xp�_v���d�5t4p���M�[�(+�����]�F?m���6y-����	�R.}�˷����(��6��zKz�� 鮂�<Pu5+�=)�ȱ���X�O�/Ͻ��8؝��67�+�s�`h����ݎ����#�Y�@��3���zt�\Ͽ�3v��_��~��[��%���@U��<%�ީՖ�衡�X���H����	$-+&��1<Z�I1 $��s�m�M"y�L}�����R	7	�_��2���+�yy����	�
8C��h0��b�?� 擲�b(̗Z��
P�YEq�!ꀂ���������G���&������,���XVAb���t�c k���H�5}��c�!�>o��@��Bep���E:��@ɿ����S��>���Q�4 �H�z2蟕�;��V�!�ד߭����B��Ձ�r��ͪ��W�@�|N�y��Xt�#P�y�J��Ϊ����D��\�#4�|t����F_T?Ot��̅�k �ߕ�)���dI���'�V� X_T|���2.@��iڎEר�����a����EK�3 �!ତ4�+�uk�Ľe8���{��֙���#��V0d� d�]�����t${Z��:���^MEU�[�8un���Xs:�Ջ��*.�Ry�"c���}3�����?`Tb�K⟦�!�҅��x's�c�RoH��.jI��,��V����iԭVA�u��n(�=.2k�2�\�:T%<� ����|������q���]�Kn
5���|uR��������!�X�Jg߳��"[�󬚽|���]Z��p#�z�.���ֻ'fe������7~�#I?�*/�0l�$I�s�G*sZ�ж|�/�mz����w�Tۍ��3�@P�*�q���|���f�h�1�_��RCR���d�ze�~��f�̣��y]I9<a�zX�][�gq28�m���FP1��5��>�W\��O����o�߮'ޏ0_Z���e�m�I8=TV�9���|��X��O��=��s�삋'������6vL����w����f�]�Y�P���e�vS�'ob���+4��u7N���uZHɡ]�� ��0XX�Ǡ���,�ʙn5}K�;,��M'|�.ZD7���l>�K��+���45���Ռ�.EU-D��!���ϟ�Ħ������h��u�<km'~��W�g�_b�r(v�uZt��歺��D��!W!Ϲ��*��ے9�W��f���G�q�!��z,�~��~�k�_�o�v�2���*x�^�Un1��\A
<p�Au�O��&�1!��]��!)�̙�s8$1�Z���˗���E!��_A��ӧx:�?,q7R����g�Cٗ�!��5�����{aR�e֢!v ��>'�:窫p\}�6�Y�$�hP���L�/�Q���r�쁬(��i���(�e݀/{[ߧ���6��2-�9�.�@�8��l6t?��TM�.?��|�yb���بݜ�'��:�e+�i���o�O^���(�h�'dP����6?�Yup����l�%�v���<��ݚF�K�}C#����0L��)؊1�ְ��2�t�!��3���n[�Rt��P����x�U���(�-�����F�Žߩ��@�.�DbT�=���R[�(b ����G�g+�� rd�A�6bʿ��#��sd[Y��p����@��^(s�ݰ���';����ӕ7i���Z&]��e����c6�L�!L�7�c.yu|�K�_
�IpO8;H�&w�RR��]u���.i@l|{��^�l�Wb�ǝ �*Jxա�=S�> ��:-�Hd|�A�пX���,���S�n�u��A���uT�"u�(&z(q�?~nz�,��|�`�⠽eXU ����w�,�x�G7������c�`Q8����|���huQ���g��i�8��o��� Ф`�ԋc6[�����&�l>C�����&�\�ͼ<rIg��qK���u���c�=U�]W�θ�������X0.���Wn�t��ݜ��(���z�����c�K��:� �������}��^�q��W�q�$�+ƽ�֨�OkM��i5��F ���g8�޼}�0��9=пZ�Cj���;i��������)-����� �$~�H�)�-tBr+ Y��̟��3��1v�0��i#�Q8���[�7��F���o�V�cA#}�����e�6�.�4E�X�� ?��1�MwD����d�O�]�^[(�����[�+����Zb$�S���q*�˽=j�(A{P۹F�v��Xi�,�c��ҡ c�f�^��ÍP�W8�im$5���2��rԄ��rY�(���A�胚Ex0�=fC�����2��¢�*�@*SD��ǴjE�Z�`��W6pV�N֫�-��~@��,y����i�U��W�4�fg|���E��a7#A�6���3��ǚ�c�u�q(��sh�F ��x����j0���5�9��|�ҵF��o��@z5x7'�� ��߀K7���[8E���S��r�%�cV����UK��s�����/��޼��r{���`��i�s�(�n
OԖןb��-e,��^
Dmp�1��؄r�j��=Ke���r6̨�wXy�%����8�9cQ+M�� a��@�����!����� MB��0�3�n@�� �������\L4���O���	� `�L#j�oO�s������1�X�clP�
�~���j�� v�x�R����oe�{���YQ�{1��-� Ye��N�O�)�F`�O,?�~�����sg�².D� 3���Qmr4p5�!5��dX�Ӥָ�F��N��%b��;��jB�h�;Z_ؽ;J5@���];ʃ�iR�5��@W�X��Z��^��j��W�c�é"j�G��9 ��2Şog�.�J����l���0)�P�r- Q���X���XH櫿?���&��P�V�RV�4fz�>KY[Y�Pbݺ�"�Ŷ��"�|e�8��o��
x2��
~H�4�!3k��ӣ�Ig��c���.̽�-Z
Ar`k����OB��-Ɨ�����c��f�3~�̻���(�墱�k:Q������&
+.:�?���-C�CGD�7�1Q�7]�Ӿ`���m�h�$a���Z*�xr.�d��
�|r�O��̸�tb�������:w�[p~ ��|�	������B�n��R���F��?�,M�حE/���|�h�7��A�e��٭�_�Q�#6�{�+���D�}��l:&�_8M����� ��y�}enڃFY �liU�~q��򩧫O߈;��r������Kο�pC��kL_V���Ő�8�p�3�3a�gZ�g����4����y�:Y�U%�E�7]{�ia�5E�c��y�_Z��D��w�ȳ�@�|�^���Z�M���S^�h�ݥ�|%�����c{E�S�_�[^RC ��(�,h@j8�����5��X�g�' P���qʓ�˞���Q� ��Tw��\�N�%K���~�E�6��c� �.��{������j*�G&ت ج�����d���1S9ț+��9e*�9<�.�,�N�ݥ���+;o��(��e�|r�y�L&v=g�f顆��]�-K(ڂ�*S��SB����}?�1�
`�z���bI��R�!ȑ��8q�HX285�SC;KV8�%`�9���qdl����5���J��+`�M=ʳ��/������=�Fˏ�����%�<	�*2���x���[��b����O*:	�C����m�%�4![�;����-�0Xt��P�iE�4[
H����L�}�{,��~�!n�5(�җ���aO���Г����$�
�!;��U�\��e�N`���Z���'� ���:�,�!�zNw�_��<��>&X�:> �;�4�N��}>��~��Is_���/|t�1��{�<��W��p�*������vtk,t�x���]�c�f�;��y��1O��@�'��-�8���-c����*�oG��4���M
���>FЇ�� �K�h ��a��%���7r,BZ�K}~0 ��z�$0?��q�_ve�94Z��X����+�^�	���3rB��z��;n�V˼���'f�&�&�m�����3K�7�i6�ԝ����������h��,�LY�w��dA���N:Qg?�`2O$�H����M���A��N����0��:���g�P��V-��6��i�u�0�����T.�AǗbHf�{�a&��Џ5��kӋ_z�%: Ё�������}Q違1��˳���d�p&n���(�<3����B����gԯ��՘�Eۣ��O&z�M�4����f�p&c�dcy]�T0Vy��!@i�MF_�Ͱ!�2	*Y���+΃V>�F0����'�5��:Fa����5�7z|v��B0ܩ��7���6�X�=զ���F� `h��o�T�[�(�~m~�L�߳=��;`<�\%E���-@� U�(�O@C��~��S�?�`�B��??6R3��6 �;���$Ւ�߶u>*���W�k���S��ZD�c��:��"*�SUI5��)m���3O ��;��AR��װsz���1 �T���K�C=��9Mb�ƅ���|=�c�;��y�{5�<�~v�/�� ��O������@���n����3� 3�
D�o�}	�0p]@]o}c�1$��Έ	�򠁜gҕ�
���X�j�s�5�H��e�s�Y����`���r1:���m���:��������'p0Oa�ߕw+ ��_���C�#_amZ�6������쵹I��~��اiȶ�
 �\�*o��g�[w�Z�9�,���_XII�B��l�T$���JnLZ��rꡣ8R�d��:�[� ��a���Pf� ձ��_4�$�<`֬:�aC[,cqp?g��p�Ij��}�SC0��Q_����z�� �������>���N�n�/���?���%��W��/��|!VT!VH���½p�s�F W6�����x�/ڋ�����
_��Tg~��,�w�Mx$���3��<��Q�k������8i?$Kʱt^�`�;cM���1� ��P�bS����W�)`�l����1T� W�f]T�1���@�m��x�g�5����U�(T�g z(�/z����X�Z��B=e=ق�D�z����S/�2n�j3��YM �yβn�ڹ�C��t�(z��	ڝ_�mcX~��Ƽ��-�@ka������&���ԇbG�������6��X%i}G�q��D6+I�s��H|�z��H�ʃ
?�_
��	�1� �^�v'wn6Ⱥ�ȯ�����
�� ڳb�AI�Nz�/������?Agx���40�UI�d�z���Q�XzȨL��X�:����=�Ҩ� pe�t���� �{���`����<��4��:�[7�)�����9�XhcWYQ8L�l ~�K�������$u����6���A�o>�K�� j��7(X�*�7�cUy�pz$ik�~��h�U_��T����~B����{D2 ��+ޛj��= �lNwmv�J���9��Qu�Q��e�	�eDjw����w�-�;6�+�Yk�u�0"<�I�D>`����rF~M���C)u��,���]u���<��[
����R2�L�U_��j�i�~gbp�e|��Y�]�֝`6|K6��/��A�TT��y��,n��
���|� P�.)α����/��Oy��l��`#�`#cP��׏�5t#�`τ^��p�_4m���[^f�Μ�i�i{�wC�>����&&�u�gI��?�J#���nݸmn�%T�@��s������H����Ot{w���<�OO �������&H!�=�˸}e��g.f�æ{4�����>��(�B�D}�����[��9�P7d�X y���/���
+��~냖� ��I����A�e����]̝����0���s�[�3u��У�B_n�]_d����R�l��,D��A�1zQ�9�\\7��cqN�<�O�ap�o�����_�ǻ���g*.�,Ԉ;Ŋ�| �𾈑�^�P��)]��g������Z��6su2.����i���DocK
�(��}��.�� �����@���^+e�o{G^��WaVfC�e^��i
-L!Hhv2lp��r�@>+��(2�I����!����-�!ӡ�I˩��L�Za������h��\�}�sW),֪A��Ș��-<�bR���U�)v�G�hw=s�]��Wt�T������A�~��Tť5���%�Hk��-�<���D��p�
2#�C�l@�5�J}v�z\�@�íY���kP>�����W�����}�v��3z������	0�"�<�"���i&R���ޔ��[&5RAeZ����;�9u	7��9�GF�[�P>+>A�-��sR�5"�_���PuO®Wo[�+]��;e��J�%!ƭ����ҵ�4�����"_���H	�������*�OL����^��&��x�<o�1u�/��}6��9����Ow��52�?���[��jc\<g�c��T )VG�J�B��~i+�ֻ3��{z��3�,��� �(u�Y�-�����F�wN�K�l�Q�m���H��ڂ���
���`���B�+O�Z�y��M��5�(c�D&���5S�t��CX�ӵz�þ�L���\���Y�26�S+M���uܰn�m�'��Xt{�����7��V6���:�Ţ���neo�����,��/j���ک}���>c[�ݴ�}�mE7v��'V��E��߹��*]8s�yI���]8����LsFS`zN� ��mWĐ��4|u�u�J�;�����-r�I�����CF<Y�qqN:���`��Q&~�)��-�k��h؄���I���yv��aL��T#�wh��ja������fY��C�>�)�XL�u���{A���:SA��ݖ��敜�=�;o{¯d�ߒs�]�kF~>������Mm��L'�3����,�:^�ZvU�5���-����PE
F9�-��|H���i�]���.��A�$�*�ete_EEt[<D�Yi
#]��}�	���T��}|LS�V3�ON�O�e9)˂���3��=hv';G�}J�imΝ\�<8J��]�~7��Ott��ʉ`W���I���g��Ԛ3v���ݳ��=F����AyH�ͺJ���_�tPqw���[��x%FȌ��aWG����:��?|{���ǉKrI0�����?��Xfv��
ל�K����v��<&�9�c2�0��M�17��	q�5o��$ i����x(���V�X��TS�1�퀟-��y�鋖��^��PI4C_�]���S�����Y���I�ia�gn�5%R��{�Xf~>�	�g74�~LMy��ven����V��� S%_4���)O�j�r
�Wv3�H��c-�����Z~D�{x������N"�6��OM�`��l��I�e��">���I|�՜�}_�y����s�f�nc-iTQ�w�T��U@�2l7m~��U�SA��5l��=��7x̬���Ύ�	c��G_Alș����A,{������Э:���|�Q�K׹C�]	���X ������ph�J�= ����Y�'�7��`�A���L�>Sģaj�����d*()y��Y�X�ucn��|�־��9���K|���N��.���{��4!lm�')��K�r��4�.�j�oi�!/����}G��Z��IG�q�_�x�M�*�/�#@��R��M��ח8��_(_f鎛���#Տ��4ݰӁ�@�*<-�+9z&�N�D0�0[=���ЁCY��s�oMenb݀䜓.����Ǻ%Q�ĥM��$���H�:J@(a-��D�ʺ�� ����ݢp�z��dVs�bhO�{���x��r;����z��}n��Y��ݕ���霫��b:��k����&���8og�������~���z6d�?,!��t�� 5�*���*��X�=$�a��c��O?����)��W� Nz��|���[*�kf��ao]wAڟ����hW�w��4G��ץ����������Mi��x�4t��Ȫ��a�Ks)�����ebG'�:U�_�ퟗ�*_���n?��u1��Y����[s��=��d��e��GG
�뺃2ޒ>�l�M/WE�����q ��uͷbt�<񝉉2�^w�V٩��I�E����'��S��� �M�x���_v=<�EK�����_�O��P���_#�|�=}k���]C�7���ux�S��g����S�M�x8x>ms�%4��F���k*��Y4�}��H�AP�v��O��v��~F0�(��3�{e��7��m��f��wW��'ؑ�`�!Jn�gzI���2� �Ybcz��W�|A�х�4��=�����
cH�.�?X�n���!��ۻ���Y�tٺxж38W�C�R�uKhI����x��uKe����o+�z&�3��� �+HďI]��D^�PR��[�� oP���٦^�0I���<-�]��������-8�3�`��� g2��Ot���/�#�(����x�Ľ_F\�wFʳ\����Nl�1N�s%������V�"�r�n=V�{���{�Xw0��X��T�b*������|��EN�_�A�D�?녰|]Qz*>����'?���]�:G@����7y��6C�����a=4Cv��Tj�?k��y41�?;܋���m��<�ޱ��}zc�Q+g���{�Y������|�����B����W���a��@�Y#�_¢����0�r�dAh��i�����C��Hr$�~��DHJ��S����	qA�	�Y�8Wc��Q�,|��y٠Ox�7	�����:vnB��s73J��7��pZ2JM
ċ����3��*��NH�2?ϵwZ�³묓��!XE�7c��1���\{X��,�'QC���8&ޮk�;�z4 x.3fw�&vK��4����86�0�Yҥ�)�0�	������_��ڋa��ǟx�1&��G��	�\��0k���#nq������׵�ʵ�գS4��˗���g�'[7k��8�XF�B�7��G������i/�P�ƪ7zE�j�X�7�_ �d�[=�����&��J�^P�(k6'������ņv+A�OH�Z��C����i��<"g��R��v�SO�WRQ���&6�.t֞��I<5�O�X3<��h�-���Pǉ��4���;K�Ӻ��U�����cSk~e9�����H���AI�B�E��]$�VU��[���������Uż����y1�)=�m�����ݳm�j<��<5�2M�?<�� ���7�ߢFrϓ[����(�'�җ�q�ߦ �A�뺆jQ(pΈު*{8q;��H�^��$�:�q>���8v�sJL���
ZxW��?�[��H��@��f?���NB�T��+ƛdP�
 �d@�����{G��P�)؞�f�z�u��?_k��t��o��6x��P �v��,��ފԇC=�����)��RB�r��P��G�.��Kś吞��{è
��ph�v�f�O�\����@�*�g��c���`�4 ���]+�3pi\�#TW�[�w&_�� �5��H��؇x�=�H��;DiM%Ep��l�b��4�3u���w؍�j�سН~�]/:��:�t�ǒ&u�>Φ�NR��T���c{�\�?��	f>�D������jΚ����CB*��D��M����|Q|���.�'��'��ӤQ�m�)q�����G��l��'�UJΗ՜4�tu�h(^b{�����|�J�@��B�j����ZW�oZ �<J��O�z�<#����;����;
b�CI4�F@��t/O`��ˣ<]�Pah��r%�t�qA��Drz_0LP7.����u�ۺ����ӣl�@{ʚHmw�6m�����yS\��:��:3��v��b���}i�dѯ8��)7T�3�v�!y:j��"voZ�l>��^3�?�W��c�J�^$�D\[�{�ך��t���Ї��d��8m�ݳ�J�mn��1���%�����w|]y:EN��Hn�p�W�������4'��?rO��vCW��ݕ��E�8T���g����T�3����y5�?7�94��iݘ���L��*׮��x9x�ux��S�9��R��F��(����CD}
��2J(��*��,��Qq9�,���&�a��G�|*%N�+�P��s��;��EŗD��L�IW������"��o`�u��U��!p<�zn[
 ��
�~�I1�\*�?�f	��H�f-�`��ܞ\��i��T<>w����c~��hK�q(�Q�BS��_���5`��z�,��~�]`��%c�,M>��:lb�y�X!����V��@��r;�V3)� ��&����?�����ުM��� �5pRԡ �X|��B%�e6�]�d^�'9=�R7_ޜ��ѫ��y,�OY�\4]s*���] ���ksR:�k��e�b[v=7��)K�$)(؎,�;ׂ��+JA�P|wZcg/4b����T:?z��O;ֳ#̊N��S7{t�zrm��Ә1q��tu,a#��VPܑz���C>�zn��@���} Y��˛��f��R�J2�yֵzXc���7�
�c("�A��p������ƽ��<<4�LXq~5��j-� �g�)5�m��8���L��k�C��x5�K
�'�C� T�v�=c�^>�����=��`}=7�%�a-�#,��bR�epJ�%�^�-_K�����
'#�v�������_�Òk4Yб�t�ܒSCJ$!��u�mAA�������(��r/��k=EA,dWg+��Ȱ��8�wv��s��-�#�a��ypw��O�>}�74��$���5���j�!�Ҕ 7�'�����Z���w���l��t���������U�qQ97� O���(n���𶒢WP��{��"膔��9���8��5��y}~5�W�ihB%�����G4��@u�j�0���z�r_�lѫ+��ܗ"�����m�8�����<;^���E!~�f/���^�z5�:a�IA�����-\\�IH�X�{h�_���z�h����[a�PU!�|/�3[�̝��oN��27��c��qx}}����2�B�7%�ޞ؀�$�t,C����]��q��n�5Յ6�,��������F�2��ſ�^͢�`%�_�B�����),���L�S�~]N����(p�t�^l ��k�B�R]�9�Q�ڇ�kk�_����q��ރ���駰�D�ŏ�ɜ���C5����o@0�$����z�X�4����cn!��R�lrjj�R��E=�Sq�$g��\��5\�Ƴ���7$�~1I~'\k{#A�kA�?�z�9S���#{{��4��p�vYq�A�w�1dQ��oN~�����a���\�>K���+)�����F;�>ˏ�joX��A�T>F����ܙn����2sTP��)¥�7��x�Gd��'){{�qb5���DD+��s�g3ܩ�\�j4�����~�삷���VZV步����_��]�����Є�C�3�J:�ZXוb/�'�B�i��t�ae�]w��l,�? �԰��J���4�Hl����[?�%.P�uy��G����9�s����y��*�a��:��){{�I��{RF,]ȷ/`�Fս �oC7�B�{�X]�sR���m��nt���Q(.QI�*+��g�]�nW��_�kء����50�����B\����7@�:���U'��1/��Ć4U�p'	`'{��f�,
pw}�p"T��[W�Ռ�_��
e�u��dv��\�.,�q�R\��u�j
'��!�:�R�4Z�ȁd��xp�I���p�s��咏�[���^��C�+����Ce�U��/E5��۟�B%�q���i�_*Ƌ�`�2�������#�T��Ri8"g=�ק{��FjO]k���J�{�-�o
�YY�)Ӻ�M���!���uh	�Yw�w�R�
�%ǋ���z��0���$B�V�{��������P�I��
������3C#��(J4�L �~��E��S\l'��t5E���݃a���p��h.Lu����M����P�7�^uDI��؟�Ǩ�� ]��l�6��.,l*���<�R[��*Q��FC�����=�"��m�;�.�#x ���P� s�۫�~U/��d�sZ�@�9b������Ъ\Be!�/�E�j��@F�Y
bG�G U���6�Oſ�Z�z#�я�La��S���e5���Ԓ��!?x��g���-�1��9�dhC��9�G(˥[6WS�<<�PO�ԲC�P�_�Ws<�G���/������D$B	Ov
YK�Ȟ��eߗ�����IO��I�o)����!4c�:�|�{���������>���y�׹���w��[����������;A��$h�B4����tsB�߲�̧�gZ]�h��������<��d)���Mh����;� ��k�>�����L����oϛ�m@�Ʈ��À5 F ���Է���S�4oR��D�����s�����&3?_�~�<i�Zd�d����&�%�E�b�n���2iD޷x��. ���k��q���۷N��%��ѭ��ss̓�z��Ɓ��<��,�v����o�k��5�ZPj+�IZ�r%�����ٿ���n(<r���G0���B$����x�ld���4�r��%�����������Y-����m��M@#�m}}�g��G��bmu���Z(({������k0_�HCn���C�g�5�&�>qk�S�����vv�2��\wr����ٜ�2��uX^��]����U�����x�����j���	h	��__��?;�I2ˈ�ό虔h���A/�n�ĭ�'�mssA��,B��G����x�m��E� 3x'w��D�5��וLb���`��c�D��� �;
��p�ϟĽ�k�]s͗#@����{�qS�G>�~f�σ�"�3a��io؁R4n�3q�x��N ���O�{������iw��s���t�͟S�t������rD��ȱ錄�����Ԍ,�W?��Z2� 朏8>1��۬���r�_��>V�k�3d*�k�'��߶m�)7�e���%���#�Ǻ>Ǟ�y����I���'��tR���	ٔ��R3����B3v�Ԝ $Q�	NNW�У���[�-/-5S��U�6��)s������תƺ6h�Q"hɺ	�6����Fo�\����	�5�:Oh�04R��8⬉3)߷>�D��\��c��)0���W�-�>8�zY{���Ұ|=ߺ�����_��V�=�����Z��UHA2�q̀���(��3�v�'o���6�=�R�V�d����Fp�eGh�F0b����%j~ V�B9��{^�@�*��"�vj��K�G}V��Au�(m��G5.��}���/��!#��.Tj�P�EeJ
�KG�<ƯDd�G�]Cb\7 ֕�,JHX�K`����9ڈ|C{����ÐO�;Mc�'Ҷ����\��i+ȣ���q�Abx>-b�Ǘ�d�70#C�`��	Bs[�O�yxd$0�41����F�/�4���n-��]A�	��X�WD�,�� {<�9�FH��.��-d�<��H�i| �s܁&tS^�&���H��cQ�	�?(�	��RoT�</W�XJc�"���M�H��&��Pu�;����WA5��	��oej3P�E&�^��0{�[�U�N�K�'a��nGD� �% <I���?��_b��p2jl��^/��K����sZڑ;��I@_o����x1�h�ޞ��FO0Ϫ��--�o'�
�����'�+D�pqb�Т�..
4�
��MH�T0�V�^�K��?KK��*���lM��,�%�`b%�=���ڍZ5(7���m�О9��P�ƍv�#f!������g���N���%���l���p���FM��0��>� ����o�t`�y�߫{�>��*{��m��@��� `�U"�{D����-<��n���3�Zg�h��8��f��J7p���<�n��Jɛ7���-�@����_�M��-P���px�����#	�@�d��11-��G@��|��Ex5���@+Aˡ{i�0����(�8F̗����˜kk����2ww�\��	5Dہ���������%�f�`�� �jڠ��ۢ��F_tzz�2�a�:�C-Ƌ��O�>]�f7��?Uu�_.4��d��E�Z�SPY`�N�^��I��Y��
�����Wϭ�[]�Ե��!�D�S~��e��֕��&/��T�P7�U���t7�+�ra���P��4�5�8O�u��hnֽ&��\p��>��76���y3[��||����n9SN�����✮� �������s"���X
PZ�e�0�o >�3�^UWU���%ޑ��\V�)�6�t�UNx��QPd)=c����~��k#���}��p���o��_��<x7$+�$�m߇��x��Xҡ��ru�f���H�oB����˪�+A�=�ba������P��	�$���9W-> ?��2=�`4���>5�HEZ�������W�LY�+��j~�RX}z�b�X�F	��0-��L�d�HIPQ	:/�&w39�\���q��wL�@�hyʌ@Ӭ�V�I)u�ַ��(� �����U2��fܖ.yg[�7�8�̸Z�r`I��xUU^To�铓z6	��##��3wuL���a7���Р(4�G��Z3�J���b>����c�nqC�P/�Ƅ"3��*�b(��6X���D��ꅃ��JΊ��d^�e�U[�6�L�l$c�L�w��b���i�T���������xU����C�UU��Y8�%�[�x9+骫�+g������H
����x��*e2�`c] 7a��gh�n?'��]�>��ы �A]1r��s�#������ã�%c�e���L�]�\�k��	�A\_W�-� 9��`e�{6�,���ήO-;5$Ԝ�b��j���:}��3�?�6pE*��c�%hȤq��t@d�"}[��8���=�6�w���a%�s�������{^y�ME��G$IV�63���X�����]�Lrs��IB�≸���g�4�]�W9969`0/Y};؋���\i�%�QA
�����p�dL�ߧܼ�,���Y�Ò~��x^E}����������DW
#EO'�����<-���>1����w�I�j36X3Q)C�rӁ<]����1�}�v.U�L���J���DO��oo���
��(�W��"$f�	Wu�z�uH�1 /3�r��� �@[Q�l?�����I/�[ f�c�>�d�Z�����mb h-}�g�P��`�&�H��EZil�\�A$�hvY�3�<�t�b�}����A;�Ryv���ev�ç�����C���.�F�T�)�9%�=���N\��8��W��:C��Dw��tv����_��(�]v�V�
5.�p�+���r9V;�����:�} �OI���W!ݝ{o��f�����5���B�8��@�ي���遣|Y���J���qA,6�6j��틛��OA�$��j_p|$Ş�,���F����r����j�X�|��K|�S�,�6����w�M�����R��>�� ��w5��*!�!N���M=���l��|p����+���􆧾�E��,Y�@�����YBi]�3QI����~9�G2g�`�4ꕠt�@�KDu��\��������h��$2U\@��c���CH0��E��3�#"r�@j<�!3_Y��q{&��]��"�g���"�б�a�\���$)�	��e'����I��J��~{==ZU`N5+4t�K���_�� 9�Ԟd�~����	��"u]Z��& ���ڔ�j���I�$�1����EP�m��c�Յ�:��-; R�V��K^��t*gln��}��>�Xv�x�����_�b�AV���������N������u��fK��>��ur�EA���&葠(�q���ҋqzVm'��!i�i5A+��;8�N�W�g��ۯA!7���sx�O�>Z�:��Hۡy���q�_���u��{Ig ןIT�}H��qA�?b<E��P����U�~&������gh��9����2O�xA`t�i��=�t.�An2Uu�5�t���:�R==��} r���P��"�b����H'N��Z��4BF��̋]��K��C�f"(B(���%5�ײ����2l~�~�u�L����ϻ����-��B5�m@����������J��ttQ�8v�!aq��
��Р����s�)���t�v|�/�Iz�%�!��.a�W�gJ��:�t ����N�T�J�(XY�83��I�wM�[3���9<�xI��\�)�x@jv$�����=C�k!-ш]�6;�?�(�oh���\O��Q�ǎ��lsS��?��A%�Y�z�
 hј�Ls�)$!� ��M����mon��1^6��,�Bv�|����/���q�(������ɿ��+�I}Bx��۬uH .�D?,��#4Ck 6Ed��x�G�:/��$=&���cQ���jS�R��j��]�b� �.]���(@�뢥.]�[{�6S8&��˽n�p�#�h���R2org'�����G}�m��6Ӗ���*\����?3S�<�� �91����܅��j	��E"	���ym�����=bm��+����V�L�}�*����R

rmU<��\|p�Z����"ĺ��'�1�`�*Xҡ4��i���VQ,}-���fހE�c�c����iy@�L�oԈ���̂�D	�d�Ds����P�}!x#�+�?pn���~�\��ut/�h�ǾM��/"�� ���5�e�v��t!G�@���^B�+����.�@\a�����>�MԐ�qCC���OU&�3Yh1Ȍ�?1�sمf�p<�_�x���D��!Ŭ+q i��]�m�'W�鍘!�?�Ek6�MAT���~�8���~��A��ö��np(Aզ�?778VE��7����f�DCf�ۘ�i�2_�%c0q�R�Ǳ-�lN�<A�8A�0󢢢��� u�'���u�s�<Y��B⨈ӄ)�I[ZM�����>�숑K�d�=�,�;4_��F ?���L�9����[���=TG�6e+�@����WS�It6�����Az�\:�^��Q��Y�ʀ��>i;:Un���:r�у*+!�S����(�|HE����
�+�������������H/��pq���ez����(� fm.�������~U�̌��e��A�6c����$�}�{����r5��}���ˊ���t�>%W�����@p+7��Ƭp�밑Y�^��$�=Ӂ�)��� �3��{����v�b��FD�SdD���;/
y���<
7�����~H��T�B������T����{kOD t�~p�A����Ac;t�쟓{�뚗��I�Vk��E�*�"+�g{y��1uS%��Ǆ� �@�= ��Vh�>�����!��|�q�f�1i7,�t�.gi1�����3j�x����;�O�;=�{kޞe	���*y��M_}��(^���.�*7*�F���a�3H��q�(7P�5rD�/�n뾊Q�����ҭ���,]e��#8�ə����R�{F���V̯��׍@�!Z�_v�2p�=��0�+bϵ���P�V�P���S$���'а�Z�pe�g|�Mm>_�Y�!jHN��`2Y�/E��~�SRO^���>��
לMm�Z�I|a�-j������n�2��݃�Au/�؇	��j� v�Ji����QM�G���q�����F�T'TF�����w����}��xDO~ϫ?Ad|���jD]@�l���ܯ��,i�F�`�a(�-�F����G�gi�uKs�� g<s:�χz���M�T ʆBc����ڙV������2+��X�:������2�`���4���B̤�5������}[�=��M��$���4�(�(��Ie�D�HȆ`�nƹ��[6��b���Y�t䚂O}�?AAr�C9}���<r�N{�^�KT��4�d��u�&�Q+�'�n�+mq���TF>��N2l׬b$9��E�1�~W�l�ڭ%���^M~�:��	U�P�������@|�^�z�*��&���tv83M�+u֯�~F8��k
j�g��RV/���xس����ՖP���)M�g����_&u��u6}֢�@c��0P�c��d!1��>7K�<cJ�*��?=6�Ԃ�M��w�D1t~����".+{;1�@G"> Vn��&4���%�(�!�!�i��=�	{�a�6�y���p�J�肐��>��q���f�����X�+z�Lm�+��(�,���v��5��x('!���quT�8����r���?-�&�����#��&�GԞ\�-qJ�<h�9E}� |T�S��è3|����]¸�t	����h�~�j"�-v^I��F�¬CX=z,��^a��-ѣ��eNG�&��p�n�()�iԈ��#�Ñ>Y����3	��ۛ���IK�嗇2�!����'nfiΩ셌T�%�'�P��.>mo^c��ߎ,�����o����Ȭ������ ��};�[莪*ī]{�rI�u� �����}i��XH^$�*y���g����G��7ծ��j"ʞ�s;��zy��s�Trl�7MF��2�>*
�m�b%�u�T"���U�U��G�����3�� ��?f�]��*g��X+�,�*%���}^)���j�H�鞮�,�|6A��:fF�������|�KR߈cY�xDV\�?�P�A%�k�t$3c��2�އ:{�g;^�����⵷;-K9EC"�P��Q��-%��m
'<d�|G3'� -S�U���ڝ��Po�C���04f�'4�\��s���h�Q����Pm�a��`9�?.*���XW�N/�|(I�hKϵ()�B��Ó$�nT_��S^������Ae�����f���d^t�[��옝��ᜡA� v̬��������j�CL|'>%�ToiBz3U䏴����~�B�9'��ʝXy�p�B͎�O���}jQ��[�vLIQ�T�<�qz`��bZe1�h##�ݾT�L;��p5wrr�M�Ǜ��������$+'%ER_Ŧ>�՝-*������Jݵ+M�"dz!/�52��vWf���C{�C
�n��=�G~]�~��>�`W�T)HkU���o�5�wX�7��;�o!�#������u2����P����k��bRH'��f ��q�x��.���/�B�ն��WK�AnAi��/]�2�w��|�77G��
��'(�|�z�G��ج�k��76�s�{���l)��ɬ���hA�J��Nn#H�\�k����F�O\7��8d�L0s��$�*��� ��\f��^��?v¦2[-��(~�Og�)�tO������X�\�~�"�dD��&8����
P? ���b|�� ��=I֝V��y�l�v�3�鶷ہxq�BII_hp��JM�n��b%A����� ��I�x�	���2�K0�\�	�QTW�H�����\KUU�"V7n'mϭ�=7M���J�κ��e�QudTF��-�	%W��9�*(��֧�O���&1��f_	d��/���d��"��W���,;8��Û	�C�a	M�b3b�+8�$2�9��0�^��-W�
�	�s��t�́�\��#�^��Z
.�.Nc�An�A�L�g���,�n?�!�3�4��H���������Q�ǝ�D9�uKjk�]�M����+f0R���i�#��
H�SQ�~�uA��ghe�t
�3�j�s��g��Ig�l��S�:/T�tu��^sy#	5
3y�x�
q�ix3�ٌ�\IKgܹ�,��ʀ/(5n*���=����jo+���.
>S)l�`�)�WD��W����͜Ø�:C�W�#�M�W����rF�M�=}�ࡔ���-����[�Rf'�d%�$����M�F~[e
v���,~��#�y@NoU&7�J
�?Օ�>�9��䝮p;�y�k�I" R�ab��:E#C��}���q��
���!����ʻ�;��V��<h?ݍL���t8��:Dam jO�?��eekv�Q��å��yͲQ�}'�pJ�p����lX}������j쾿ˈ>:�h���"P�?t=Aj��p�[�]+3�k'�iWa��3<'��^̓?w�	����2 z4�K� 	#��sm��s�s�Z���nV=:�?L6�ܹK�3�l��'(����m�G^�$����C9NLЂ�]�yx����|��+�Ꙥ����{�٤O�:ҧ����U˻0�qf@n�$��OC���)�8(�O\`	��݂oF�V FI����P�㱁I����cGlA튔 (�b�E�p�8���Lyc��P�i[
yk_��$�@�ޤX�:����� �`�Z���J���.���:f&��?_��8�����W��g��b<=���Y�a_�djR�{㷪I4��abYC^�����;9�$£\�q*yok�6�r����_���ҷg]��5.���C���߃U�-�>�-m@��8�$:%��ep�!�*>3<�k_5�VB���C�J��|f��{⹫7$�v.�ٙ ���>��_~��#q���=H������,R����Y+��0�:c%%�kR���"��q&����R��V�ww]�5�K��,KD�LH�[切�e�{��&��`�ݣ5�G��|X
'P����Ư�{���@��Hd���C�R��l�HE��(�F����^��cs3��]�������E�]
Ww*�eS��r^�T������X��~��F(����>7�!���w�����Ak��O{���	����:jc9ˌ2��o��ǡU��O�9�c󺐡�k�	]���'�^^�3c��L}sL?����}v����ڙ�w��ׁ����B��<�����Vh�(�t#�	h�9�.���i���,mjT����������������e�0�����s�`^�6�u��k��.P&Z挄o(]��Xբ��h�:A��v#��v��k�h8�h��7a\y�g$!��Z~��6,R��3_N��;f;�XyGH%�
<����/��ݴ�)C�v��J3aJ�Lh�&�2�k}1SpvD�|>DJ߉X��P|���R��D��V�F���%��	ʨ�A�Y��{H::Yr��L�=��[/9�iv�ۛ0������yr���ӏd� ���K�
8: �(�.�D���z�#�J��@膦�v��}v�=9�����9�"-P�E%������<��V�$�;��ߍ -y@�.�d���XHXH������ѥ/cv����_�h_F,�B(I���Î�Z�I��,~�u�#'p�kХ�����$&�,G���cT��GB�3Kmnp�z:���<7���_]��&��'T(^M�/��k����#����u*�9�PE�����GI�F��`gCCA�ngZ� ���S?j�|��Q�K�.�Qv���g���[�g��Fu5_c걫�t""b�\Ei�:�t�킵�g9����ܐ�[t�8��}��U�>���RR�w�JO��9�x��.�EV��l�xR��m0�a��9ӵ��.z�N)@�w�cJ3���eR��<+l�:�Y�z�2�]�l)Л?�u8>��.#��g���zU3��>�MQ3r�nRi� I��W&�RgHڴf�J�� Z�������OW��Y�H
�����^���?U�	rz�U�Mq4�^M ���l>A����֛ޙv�����O��X-*���kY���Ŗ&uz��6�yA{�)wj�O3�k�!�ÍTң�>��� ����X��םi˰њ��K��Y'zJ��%� ~����o�ƛs�������r�~��t������ � �Ł���/(T\TB ��iuY�۳�����$1΁�_�F���B���L���JU�����	pHx�ZM�޽Xn�<���^��m��4�7i�/k°�� IR�1f�Y��0�?AE���������~���7fU��ɳ�-W9��7=�Q6���8	F�;��xڤ_L���&��`J��������ԓ�F_��Mv���F�S[�U��bi�T�E��0��h�A�aYQOd���@(���H+���Gg��2��5��uYY��,��˃ڒ�dj戴���b��\^�ܽN�����+?��Qk��F&ޓ�\�ذ}��"��an����(�:�O���������/xZC@"�t'V7�NqEE<-�E��O�hu^���ִ��%�z����:�]���󾑹ц�s�r�d��q7�w�DYAO��Y*~��͑l����D6D��5�՟q��M��y�p'�?�2$g�-.贅�(��=��Ͼ�z�	ݹn% 
D�g��]�����T��`�yR��R:��n�m}�_��@��!�B��Y�d��O�����L }�U%��i�)<�a�e��P��l�IՆ~��ڪH�cý�ӳ��js���H���uW���J�s�fSih�����d�'�'V�6�O:=�sѴ��Vn�gOH���S.]Q���ŵc"��\E2�!���P�D
1>T��J�	�7\QQ�tGyz�h�ط�x���IHx����D��<�8�Y;.���m��jY���o�[���Th�NF"��cSg��5� usS�ڛ:&th�cLG����$�-$ޅ��n)fҾ�1�}W�nx���u��oa3�����&Jؼ����qz���q���q��3kNNN�T���pu�ίB�>�'�$��t�zh�G���R�:�X� ����Zm�ԝI�ߢ��t�9�87����m-��CC�=Q��' �W�<c�8v�wC�-����C��]i=�!+{�E���G��PgC"���Y9k����ኃ����[1��Wĺw�����5`���Au+�����@o��UU�ɛ�roS]gZ3��(�p%:'^(yCG2;A�kT�W]���1���v��g"�ZZ��M��4G���u���O����gĭ��Bѥ�{�p����|T닢�4�'����i6�a:El�N6Vإ�~4�/b�\��}*(��朚��r�'���^�}T:;m���u�Y'�dF���Շ�A�K�k�%1zz���:����B�H�6	j�.u�8�g�/B6���<�_�	Ci�]�	yVp5y	1��$_V6Ԫ����.#-�{�r����p����b��*�7޳�)f��[������.Ǫ�t ����vA�Y=0y/OZ��YR�/q�M�u��;�ݧ�ٴ�#=c� �
(�Z�d*w���"�6}��Ɔ8���y�V���B�f]��S�jlj7J��!�c��kލ�b-B1=��(��@�t��p���n�R�´�9)Պ�����K�V������!���̀5ǰ�m�i�g7D\"���L���{��B�-����[^�����ٕ%B.�xS	�fݚg�;/K��K��6��&ZZ��A�2����&I��c�6ixkP��z��MW��2<D�E����r?���e2gj���� sQ��`J?��	�������==��G�a�'�d�1
����g�	���XHz���,�6��!LK��{��=&��3�{g~]��n���ր��޹��_��"w���hWE\��V����o�:�Zh������l8|��@
�J��P�	$�S����p�TTe.�.s�34;�Q}����-%"�����K���XB���fF���V�a5���r�lN}]4�R��5��gE�!�'�%C/͌:&g��_��x�{B�DE��5<eWh�$�-�6%��u'��V�E˝�i�ˎ_���W�j�3]K0s����D-o{��'�bz�>�N�@j\��ZB&J'��D���g�G�~���FY8j�<�)ФT�`+j�R��"ٝ9�����Ǧ=��[I6{3��;������I�l���Xj9ȝ s���ތf4�T>���?���c��I��^x�|��q:�
���� (	�W&l@3������h�,���mE��Le��K<�!?wN JL�@����t�Zg+���'p �*4c�<��-c>��O��"�[<�9��%`��h��Vn4�0Q=A�Y2����$�-_W:X���յ�{\4K���/֨.�M9$�g�G�gK�a��I���<4j{�m���a&�l�����C���p���~]q����|;i��ى&ݹ�\�i��M#�x�����~t*~<aI�B�s��5K��A���o<�%LL��%�����W�4�wD����E5��)Y�i�j��������vHl�>f��=��b\G�<�Q�e`�Emy�r{{��@妫W��G�G���"�@G�:��h�Y�"�&F�Cw�fI˥�վ��c�؃�
�;���Ƥ��M�����u�%�nyU�YA'X¦_R=�Q�E˩[5��g�b��5[�[�F?�h���=�X6�y7SR�;���I"�M����7�Ӎ����M'�xjgO,r.��s_�[cS�z݊�c�������E>V_��X����`Ե"w��c@=�loV���Pxv�خ�Ţ��-�n���	���^V���/�䓿ہ}�󳵍XD��T��ms��2�n���
���✖�If��uta��^f����`��?�^xTq����y2ZT�ΰ@��qѕ^����/�E��]�g�,�3�Y�vCٮ�Y���t�=�y�Y�qt�Iٯ�g'��&��9o����l��_T��)V�RhJ��4���n���H�L-�G)27s�ǳ:I��Y��I5?�YR�X�F��\v���;�S�m���k˽�����;9�C���7i�]���8歕)�w
	����]u�V5z��`���	BB��}j��Rô��+f�~@j���a�0�!�N�g�4Zv̤
�B1]���$,���f�����e����ە��XD@��]?�e����綪H���3x���q�/�.��)_m����͎-��yx���,�(��1s�Ǎ:+�C���K�O�Z�W$�F�*/�y�.�b�)Ø�2��f����Sa:����F?���q�G~��D��9>�t�M4�v���{���#r�	�U똩�c�ʫht�g�u1�x/����es�h4��L�?T�{tnt���v��W�%Q,��vo�N/Ifv���{f��;L��fVE���G�/��#�.����"�[b��'Zj��?R�\��_�c���U�* yKmj�|^h���L���U��I�&P��̊�}�7z!)i����Ì(���s�Z�z���7��uUڽ�o�3+ҿ�&�o��j�|×��b����V�u��#�������&D��nX���(����_�����v��jm/����LN�n�m[p�bnqzǏca�! ޅ鑹��%���������h�5��E�������$�Zw�Cَ�/�uh�qU����w�2�p�Xտ�����k�Ӳ>���3ή�t��IО����W�wwcS�,ރa`��dㅫ�j8������[˅�鞆0�R2r���Jע�x� ���x���s�+|�����a
�M��/�.z�ݢr�G�
:ť_Z��jǡ�eǼD���%k�WR�XL��f���)��e?��v�aXN�mM����-4'gM�L.���f���m�4"x�z������
�g<���vy.��E&v���{�X�o�"�
���0�SJ�]f�:3�8�[��%�6k&�9�Qa�|��kc�VK%�� M�_�0�y-7��CW�Y��)�M��w�����#*X)1���x(t�dЈlʉ�~��]���)y���Һ�3���wʷA���v��=g��[A���abڌL�F-k:��-~�Vqyy�9V05�Z>�:l�oG��Ȯ�f��h�O��=�n��S��R\���?e�;n�&>K���v��(�`IE���_���i�=��'*j��9��d�p�
��Y��.�ԯ��+�Soe�)�S����.A�>�:�p�Z�����5웳�ޡ"���έ�'-��蕷�rI U�O�{�*�������e�������+����\�v5Z[Ӟ=�My+�E�se����4ߵ$�?eEభ�1��
KI6��;C�睎��YF�=ȜBjZ�� ���~��
 �Ȫ��#̱�/�E��r8k��`G$Ѵ^(���:���TI0���F$�pa��b��]&GDd�$�x�����<�OMnw���{�^���z�sjΟ58y39�>�!22s����W`�+��b)��v?����X�a������e�������|�zVs��A���!�s�o��v\L�g�	������2 �,ƃ�l���š�����;��	����t���۞c��7Y� 'v��ΕK�R�7Qҷ�w��Z�I�<O�mɰT�M={WW��Ee��a�[�K_��b�>��y��DAH�<e��y�:�&=#��K�2��OJ��s>M�ϙ�.�x���9��P���s�#�; q�1,����KP���㷦إ�,�Ym� ��+ ����M`*6}N����԰{N�[2��;¹jtQ�f�-����}�B�[2F��V�h���2At���gl��;׍~m�Yu�+�2�	���K!W`H�[_6��EVk�Yb!���D������g��;�[��.����q9�n���(�H����B��A^�����I��=l/�D��^��h�cQM(�_ZcbQ�;���CٌOm׻�5N�'J�lm#��]�B��f	������4�`"@�#��o��8j����}�x������Y�W����,y���|�66��J{h��Y$���$�����5�� i���G�e�J�}�l�uk�4W̻�~����O�.�	�n��Aײ���F5[�z~�wo���+"8,t��e�7�_��)������}4�1�ކ�F�A<pP�,.?G�ï��?�8$z0��,u|{�|¾m�OR�^�pFb��(�G���<LM�.������L@� ��?^|d]����n�Կ�����J��1�(��B�o���QN��f����e��T���h�ҳ��E�]�0FP��Da��i	V-J��u�»�k��P�ɛcyN�Yx<Sb2�K@Y�M:�w�n�"!sse?z���l��L�0#�'��n`�� ��G�&����<�������߶&���4�h�<�̊�m��20T95��i��?OH�	�'������}C� ��h�'�s-(��p9(��gM�_@��30N2��͗F?�65GȮ�,��r��3Nb�(�V��7Zs���*�Q�U�F���ICޛs�����c*E�d�$iD�f�A��߭k��N`Ys�X��
�r(`�H)�F��Z�Z������X^^ŝ�&W�sa]Ե�p��T`�I��f�+��v6/��aR���O;bG�%�h�����`K��X��d���h?u�|���4�"�u��+yC�س,��Mx��o̝�}�Ǖ����&�0�)�$���^�ɳv�u�K���.M�D���5}�������gM���[+$��v[/���"�I��h��w]�}g���N]�w2$��@�Zu��P.:�wf3��b}@������D1	���k(QS��s{uOx���p��Դ>{�ë�n\.�����#�"3�#,Z|�i@���x`m�LJ�M�B����kتӳs���m��0X�A��l@0�aD�Į�0�~��0�[��7����Á�2S�i�&:�vmo�i�?3��(��ϹAf]��B�|��-=�dc,�� G��+�*���TJ�53M��Z�9�&B�V'�r$<��ڐo��JRe���M�F���E?O��/fћ!5��fW�������9nP*e�U��"����6;��Ђ�2U`V�Z{�i ��4��g��У�/^� �� �{J��M�y8���^��͗;�B�L��}P�5ڊ�� Ņ.�e�T�2�5ຜ��YJ� 9l��L�de=h�]�����rt��g(4�@���.���4|��ϻb
�ax !�Y]����T؞)K������K_�g6�^�G����4W�6����wA�(��#�)[���g������z�a�M���U�*ӵ�?���Q�AP��|��|�P,�m�s�Ű���'�Vj�l4� �x懟T,#��+F��L��O����^�!1,������ɲ9"Iw�O�����9����Ui��t��@���m���S��k:sOTc7*8��}��v���u�����zi����Q"o9�=4>T蕬b{V���?�ԠP�����q�O��\n2��?w��f���+�-�=����p׭ �~���
/�k��A��ݱ���2�r�ǟp^ԨK{�Sô��8�
D��fX>x�>;{��0b�r2ܡ��`\���5I+莾��������֟4=���L�E[�E'w?�V/�"}�$H�V�؊�O���l~.�a��2VӍ�s����ኗ
E KG�v݆Fge!�n̿,d�,�y��o���ꑋY��k�]S��8����&�xg�W��WCG�v�42�Z��SC�����	
ڱ�d��u�uiN^�]��L�)������ኙ1̠��u�- ��9����,̸M��bb���ݭ��[�ڹ�p�^���������rٿ"JO?�^u�!����|��G�;���.~.7�r��OR�X.*���c[��*�	���?�,�M���wB�g5���Tf���z���sv�����Vπ���H����_����.�gF\f2�.�0pz˨.�|� �z�^:f��Z (��i�E�j����!G-3x��c��9Q[���kz�<�9�Ӿ�З����,'�Gtq=J�S��c|]�����Y ���;��?|�����$��p�cL�ԅ}8Y����I�B�^@S�:(ߥ��E �k��$�۽�{�E>����B��\P��ڑ�D���g�	踄X��%�!�h�2+� ��%��s�� �X�4��ZaUl {ST�,��C����br%[��z�nG�O �[Ԧj�.<B%:�����%�t�ѭ�5K��Ǘ<3�К���,����fE�ui�����"..<9e��[c�4��u^;�ȅ�+{�[7�KH>�QLt�l��lV�+�@/@����+�F�JA����9P��Ũ�֢9�k��d�(����)��i�G�� ��G�9`�Wt~�͓Z�E���H�\��!����~�Y��*�`$���ʡLY��2��[3�u�X�,П+B&<�VG�����O�s�?�����z��1��۳g�f����wb}G�eM���kқy^X�>��Ӣf��(�\{�sy,��6vT+���v?��*)�,?W�h�^�8ُ���$ ��o��-6�2�g��%*�jo��63;Vcv�����w#h),���ؗN��Ɖ���������`�{�9��2�
������OW6H�;N�\ u�tZ�Y������)��j�%��D��u��7,�_S[@ݪ9�`�.g=��=�H��U��k��B�/̊�K���"!���@�M�� �ޛE��-�ܭvl��Z_\HcP Q��R���~�S�-�r�_��Ujm=�.n�/��'����#т��/���������nra�=��z����b�h�@7��ܕG�.Ztb.lV�\��J����܎��~$�l�b�yV�ʎ�Zb:<��~��z!���K���B��y��	��7m:Xس>Oڒw+�ж��J��w��C��E	[SS:�<T-�U�����a��>�X�G�v
�h1�����쇊�"�!k�N�g��N�>RYX�'�W���|;��`>fӯ�p�W!��R��r3���$_��Ix*�X�ey���㉢xV�ݝ��%RO�~��"�&�w��<��gV��=�D��W�/R�:��������vB�|��3���~Pn휋/�a�g�O�a�LN���m�F�)��`Y*�R�ߝ�0�:���{��#��d:*,I���_�uP�n�'�}��f��Cy���+��no+~�'r�z���1ܫ�|$q5�$D}�U���)]��;���:!H��?�^7:e�tV�9�ś&>�$�\��&�2u�4	�R���K����v�7~�ڐ�����6~o�����$�Fp�aU�q���V�i{��;S������*���!u{��[��s;��j�c�d	��f��V�&[5���:� -���ocF��,��
�����}4�K�(X�f���-(�����W��V����57+|��~�U�|3�(��q3F�Ĵ���m[�G�0A�æ�x�����p��rč��;��_:3��t��p_�tj��?�x�+1i�7G��ޔ(��եy՘��?T��#��,i���l�!A#������8��B�o���?Җ_y���X�U�����p}�?��:,��{DAE�E@�AJRQ��.II��4�G�����Jb���$�`�y��<����xyy1g���}��^k�9@�}y7;Q4%��3�\d��{��_N�^���H�B���}YeX���A[�]峐'�|�`�Q�t� ~Om��.wP~���?��אv�T� ��;dږ,rDe���>�CN�A+?�y���si�,��%��n{<�9����%� �z��|�]s4�����ǝE>��a'4�w����@�b����H/�X����w�		��w��G��-�O�CK��9������8�8f��P��G͞���y��8�o����N\���C8!p)�XZ�f�r};��w�$������z�w�R�|�~����)Hv�����"��~[GGg8�pe�G�bz6h��_��q+�mY� �HA���?{�,
nE����;.�U�yrs��9D��U��>���T�Ĥ �,,��֨炵ۺU�}c��	��[<����FW;F��Eo��k�V�����՝��J���B �q��y�|�|S�D$ dθ��^���ɣFw�ݧ#�n�ē`�.����_ 	DO���K`�ɾQ�n�U��.$�|�:>B�d'bE�y��6���� ���m�W��v8���8/��D��]�`�Z�v�ی�:�f�?�6C��Z�YN�����
Џ�s0��s�Ah��}�� ʅ�ȩڋx2�4���홓x���ס"((�����Y����KST���(�� ���)������$��'�}�-�j爇�W�8pؗ�q��FvM�ģ, +�?�"�Lz{����%�漨�]���!Ga���^�D	�WeO��Ou{a��"���*��98t��!HV�exwP�k1�޿�y�~�N��YKE�D�����{b����E0C��r.wb�;�_�z=��o+�����J D�����R��r�
ѯ�Kɔ���,Ѐ�M�,��Fx5d�O��ѯ�zH��������l����R|<�V��+x�����Q�ӧ�������..[K���	��G�Y�@cQ7��2nm�+��ϧ���c��&v�:�����{��9.-�,SM����ҫW��h-�:�N�$;�3(k�������e��*�?�j��WZ7��(uHT�^��P����)�i������э�*=���K��/�rfڢ*���`uwO��)�7q�svW�'w�"'�9�DbwP��5Qk*���%*�$V��l��)f;��9{Jٳb��N�c&���,���I7�+��4s��p�b�cwm��E������)R�YςkJ��w���R�0��Ώֈ�xy]�C�@Z{ըw4n�7�����{����>���xS P8�}/"��wB6=ȇ�2�� )9��e:<����n�?C��\a�)w��� b�x��X���+���C��}��.����h����dw�;̡�F�����v��c��>��Κ�+��T��2�_5Y�:jE������Zj;�Alnr)�^x������[2{}r^e�[���1y��^�%�D#1��p���'�4��o��NI),�I����iHx�̸����6H���2�"���>���c��=S�����j��eW����e��0K.���"�:Wٓ�M���J,���1V�8�l��:�<4�@S`���s7���ZNlPKK��5�3;��!����g��ޗ_l-W�	��e�-�Dॖ�N6,��o|{���d�<�"���k��@r�����ƁCbخ��|�T1&��UN�7T%�Zak��VX�BBO�1��3�x��'����Y b\�@3�()鮑e�����N�Q��Z
��(��jCYWp�R�Oi�����;u�[�	[��$�K����$px:SH^��
U�Jt��{ �@2�Z�Y��3k�~JH��H�_h*#��xm��)���&�7���f����V$�U�
xl��y���WM��+=C��+�����ѸO��cw%��0GNw݀`�w|���|quS��`�'5�E���]vW��ĩ�	�K��̉IT���e��w,O`��,cG�����xKH;�x�W~]����P�}8����p����C�~o^�vnع���5
��2�Z�=ѵ��v����>��}v�1�L����q����sj�!.mΫM���/�S�J�����{U��0Z��g2ҙ�$jf%P/�%VP���O��8+��w��L�MX���8��w�A����aQ������5�C}�wJ����CTbי( �m�����Y�%��e��r���;��F3�$��EA�-�/�E7N@���&�]M(�C�E�"j�X�#��_Q�׆�x�"73Q>�%	���Z9�����sG���Y�1�9�wx�-���w<���-XOXVơa?�w�
1�e��+VA�49O{�#~�J�b�	��>�1��ןg*�������@��g]_�����L`��֔N���(�(�*�'�i<�3?�<�bp�EII��.>I��3���l5S��	œތQ���[fD}U�f��x/|Z�<ۢH�쇈�v�����\WU�2���qy'_Ֆ�Q�O#ݼTf�h;��a&A�x��Z�е�_�W<��h��]�7��&,�o�-�.��g]AA���ݼ��),�m��9c2�9������lP�f�I�y�w+�d�zr����0㗞������=�����Ft$��R�/�DC����Ą���7��jj;�����~g����xcj�7,��r>Np���9ahdc9 k���^xچb{n�c�O䔂N��	�p�ݨ�:bG�MA�bR&�B︗�[�5:�/�)�\�d*Y�'�{`�:F?8��S�P�e��V��V��\/�]#Ǣ�>����/���_��-�bf�����7�"R�I;]����Q
~c2��;���)�t��J�B��]bV��.�(|��<e��2fw�T8b/39� g�Aby��E�a�u\�2v9}8�8�����~��FY5�h�0�w Ȩ��+�A���51���J��ϓt�Z�;p�P_��b"��j���?�1���/��2����:9u����U�?]5��YTFu�mq���x�[��~^Z���X�����J�M�Z��]A��ԲL��5F4���Y��W5�!cq�,rq^�>�������3K�A�χ�jČO�u�\f����t�ݘ�Z�����>���QSY��W���N��գ�Cp!���dC��� *M
�X�P���XeKdP?Z��1P��CQ\�zG�lN���
~�ʯ˧�&�-��=)�m��%� �An=��������˲�w8Me	�����Hs+�o�V��*´�486ۀ70v}��g;fџq�Ӱ����f�)Gwj�`�խz��8R�gh>}S�KC�g�</d�
;S�����䯏��e+��'"��R�����,�e�bK�v�-PU���:�I���V�i���i��n� ���J��K�}�����\O��9�Y�^8l=`|&���_%�]��j��v�\�o�s�F#&�����0�g��@�����}=��w`�R�S�p��� ����?b��Io�])���Z�N�׊���`���sr��}
'yg�;�ٸ�\ʅ�.�
{W�Ϫx�H��07�v��%G�w����]��@"�R���+6�S4���\�<X��<PռB��N�TV�Jp�$�$=�P_?�q�9mɷ�N��}�����q$`.����un�}UG$�sGSՠ7O��A$y+^�K���\�~�|K��_��9��>M�:{���͂Ad��M��2O����Y\�������5�$��АW�/K���w�J��3��{�l��*4A{�|����^fS\��ɳuȬD��&���0��^����Y���M�	�Zf�������,g
Ҹid�;u,��'M~�p\a���D��v�!��k�X�9j'����D||Ӎ��x���Sq\�1G4�尠�Gʘq�mX�q�Cx�+�s֨�^lR�<3��Ь�<Eqݝ���҆�~U
g��]k$+�#p�o��=ӼW�&�R5va�!/򉰌C&�↯������B�~�ă��;�`0����GyEu�
��6�`Wt�2���Ts�6�v'��=����ә@�"c�w��쌺Ys*%�)A�L���!�7�0b�z��-�-2x���W���Xe�0ԉ�Ɉc�}��z?���G}w%%
{��/R�A��9� %:��j�����M��g��Q\)R�Mb�ų�]�aY�qT!��Ƅ�2<"W
q����%�WM����8��j�8��UvÛ�DA���*/���	�XA�홣h�z��Ԟ5n����ƔI��ry��<�i .μ�|���}֫0 ��I(���!b�<s����J��`���(�ӿ>U}a<j+1�s$$��#��Ӻ,4��߅}�[аע}��f�`��s}�6��;��M�3��$<�Б >�OQ_�y�Zԏl{��{�z�����
��9}9v��%+M$���p���E/����N��N��kL�C��H�Гn<cX�\���/�L�����O�Y8�pA�X�wp��~H-���\����pض,q�/'A�:�����V��5��:O�u�vG��8b�綦6{����R���w5I��<����l�j�ɧg�R��P~8����V����/e��t���w3p5u�@�g�ӡ�9�@,{��>.�I�����;{����"�Z�?��/s��@('���K�h �8w�K��)�-�`�uw8���"^	e[%~�W���q�(��\i�	�J�L}O�34�oPk{�;oࢴ��zN���We-����Т��S���%�¡�{)΅�ӧ�45�֩�҇�@��'�����]0�{-f}���>�:��}y��5i3�<O����a���rx:0���w׏��D���I��<�o��-��ځ*�lo��0����� ijz}��(�R�ng��d����$f�(���浑gf���;ļ��	+1�_=X��8Jb~���/Sf+Z��-z%�(�~,��ܓ�n��V��y��N�:�"���K����vW�C86#ޜ�a����`d��f�o̵��X34�g�JM��<�=1:��<��'"��jC��.����6�;[kyu���A5T�&�f��3K�$�:�<���~ؓ�a����F0�v�����)��~K�SV]k��@��s�: �'��qB�L��R�)�eII���נ�vKbȏ3!Rqhqw��sU��^����ZyI�\�k��,w���s}�v��5^ޛ+�Z}��q$
l�FL�U������
�sP�5w� �@ �fd��Uc��0O�/���Yh`�1����b'�n���=Ą�_2ߎ.�ogbFy���k��k����F�p+U��qy��m��m5v�=[S.U�%w���g�4��㋪v�P���}V����A��l��y��q|�}� �~����)fq�&)��?bbV��H�)*�v�	$Qp�yRC�k>,��q�ȴ�CnH�t�D�袡-�ӫ�Wi=�3U��$<}�'�J7dO��s:����T��j��� ����>81+����i��S\O6�;�BBE���3��g�C��ߒ����։<�{M%���*�@���O�6�E��|�Xp�z�i��4��x^��T���43ZZs1�}lD�>�K��~#��)�%v)�W�j�㇘`�
�TX���1�c����G���}wR��wܷ���ǄF�ϷX����r	l�8Ծ���78`�A�柚�i\�,wAW�vKH��M���͐��B}�.v�c�ԙ��7�+_����s��@�=	n=�d ����.y�V$�ׯ:�S�L���=6�N+Z�A�󘔔%���%[ِ��ND�,�(��f^���bgC�}|��W�<<$@>>�sU�Z�A�z���F��c-9�9d��m~g�^������Ξ���e6�s��}��0��EF�Y%�a*�� Y̛�{�rE-sn�{J+EI���k�AH��&�F(8�Dr�I�YX��ry��h_��k|5�ס����ָv�_��9̲̔?ix��]w��Ꮾ��K�^�A�ё�l���b�ui�'}�c�ʲ�������,y��A��������w`\�<`ld�G���NJA���7B�5^����Cc��([�޷�458}����:)-k��`��qGb]8�ɻ�2�6�5��
u��]�|�-T9M�w�m����^mT�ij�L.w��W}=��(3�@�X&k�hZ�Ϳk�og��4))(�(>`�&�z��Vj>C�x��~؛�5�a��\�d=/
2=�ʳ��ۆu9gS��\��R�z<�3ē0:{K����R��X�e�$
��>��Ii��b��X�_�0���Jӛ��{25##ug��4=�?:�XgG|�Av�kp�Khjn)�/�/������D��*Z��F��H3+��6�^��]�ޢ��%{u�%�l�%myM��c��K�h����w�C�����^�m��r�I|q��f�7�
�r�~F���;wB)|6z��-`KfS��õ��ʒy�n+s�����.^QZd��춓E�Y��WT��G�h��r\z��h�_1
@A-��އSW�\/ }������	2_�e�Tfi����n2���v�b)�Îu;u��.����r��v���Aibۻ�=�t�}�P���ۯU�K'�|m�)�:n�q�ʬi��Q�P3��R�I�7o����E��a��-���2VG�������q�)3��$��F�b���J��5̐��UTvTV8�Ȟ�:8���П��7��=�|�C�տK�,���X�k%��5�X\Y�y��;uqN۞��Sx&�+p��o��Lo�0lMLJ�` �ԘvǑ����`H�_�ў�f(ΰ���#��x�ksV>$d�ͽ㞰��JQV��#Z6�C_T_�|�  �T:H'mpl�m�]��u���Qѕ���C=�g�6����}�3i߻Uֽ� ��^�w�d��B����$��x\^���v4��26��_;qfk1��ˇ�7��W��t���,�gZ���ΕTf$�r�V8�ĔHoo@�/�-]�FS$1���#��.�a�/N-t���ר�_gnn����`1�{XB�{�H��cԡɤ6��
z�e`Э�bt���4|�#>��&��M��ZR���#�$5��Z���YB���A���b�7d!��^P����pe�`��m`o���ߊ��;Il��N���Գ�����ڗ���öRQ
�^x*���fb=���Ԝd@JT��	��#A��c�as�X��QzWG��v%���z��d��U�ڟh�H�|��h�M:�L[V������_珗{�o}+���BL�YS�_�̙��.�F�!S����N\���@,FD��K��{e%�&+�be�q�[��2mS��Qx:�)��Y"�@�D��k���-[�|�"�C����4��C�AC�)�[��<Ej���������	�,22[n|�
���)��[*/ {��O��MA�pm�e-��q[b1w�z��P��k����!�y�^[JZ�&e�l84`$�@����|z�~N�IH���.�w:�Ƃ
�;��JA'��ꩃ\���)���"g��<�ge�x�&�ֽ��&�D&�./��o�6��E^������gM�8���hA*��Q���͑r.�G�6b*	�
�X�$b�RC�<��#��B�W�]��N .T����xM��fߦ�c��J�:V���:띞���M��(�$�m�C�^�{Bi�I���>��q���7oj��*�;�vwo��^�h���6���v�Pt:��x��1��W���AQ�b�@�[n�C�^M���Ҿjj�4��d����^u�6:�8�E4+�����N��Ó/G�1�gUC�bbp?�e8��R��~�J����#�T�sv���Af�Hsy�{�>��Z���������}���o�[O�{�Bng�@��ᔡ߅q����?ȉY�+��B{3�����7J2?ɚz�����M�>r���׫̭���U���RD��kl�˭��'�XU�UWΫv+x|~$)�VOl9��R��Sw[��]�S �Z��XϥãI��n���"�;�U�P{�
'' ��M$��7_`�(�Փ��M/�;3%�eq�c����}x��j�A��p��ҏ��X���م�R0����P��.y��w!ZL�\�9IM�#M٫�7y���\�����N��YZpK\�����4%Z��>"�DrI�|yW�� �i�a�ŶNV��;:���է�
�a8Vi'b�QY�^Y���(I���lLW�9z�X�Ծ��r�ۣ��3xѴBP���JK��+f���5]�c�v�ݑ�]���W�F����R�X�%�0"�M:)vv�����#"�6��*vm���N�����ط�x|x�>�W��싦����/���9�+�����g<e�8ȂG��,��	����X!l������� �e�ݜ.a��NQe��s�����6&e�u� ;����A�{>�� H�=�֧������K�A��-#b0\';}��g�8<������p�*�;��O_��kW�K� ���7=r}N�EM��51��L��NYD�<+�|�.� ��V�J���>��0�:���R��1��ۓle��X���hkda�b|T��[�Pw�M�?�������xqj� B�cH�/ՠR��ZsߌYR�g,�斖�������ɑ�#����J.��҅w��
�����֞nJW�u��\׽�(A���½pF=G$#��D�����.Wt)[�aW
w�~��(ߜx����{T_iڮT؎�_�y���J�F�����|C����Q+}��
�ز}v��<��[�KK1�4}rvI���cC{��O�dq�C�>�h������V�xEݘ�|������#���('�P%�`WEUo2�p��Q�䴍U�/N:Npb�@�
sԻʭ���4��	��&/ ������ߋ��������t7��$��(G���W7��yH��x#�q"pKe"�%��'j5_��ks�'���D<6	}L�:.`�GP��5��.JJy@C��ᖤ�O����� �<5#�ظ�k�Z��5��Z���2[���d�DWyW�U���;�;QR���x��^�`�(�l��^��d�ڟ%���Y�@��რ˴��@Ա�Y�ch�tJ�x�R�R7zrjs������u���K��q�N�\i۱nq�S�(a�d�i]���4��Cv�?ޮY��bd8�L
Q����Ȃ�Ȯ������_%�ϝ�/�Q�\f��{�
�U��՞*y��f��a�6�@F%������U�D1os�+���R��E=��{�G9���+�lA5�z�ѱ�D���)Xtl�+xCQ�h|؝̹>f�Ha�O`��(/��Zg�66GZ%�&���~��
M`
Bed�b����MΔ�a����`qA �g+*�-�ndx�_~�����.3e���;o�������k2����p�	��>�2P�9V)�����-	��O,������Sz��i}�P|���ze��[wY4��mg7�C(�J���{�3�- C(a@qʫg�����;���3�V�N�*����Z���_tn�^e��'��~�����@ӥ"����ROv���Mi�g��#�����
jNO�����l�����b���7" AB����m����P0�(1|ېK��Rc{���a?�kܙ��t�_7�_5.�'���"�1!>>Z�N��"����G���+�<�[v���
��.����ևd]����+���	�Y~Xz�F|��S�Y���;�k�]45�qC�O��a3Ϗxy����dd��t��Ź�����L������ԅ|Gu����B'6W��.��j���t��h�i��a�U�����r��McuMs
u- jt����Ԍ�x@�y_'��;��YM0OO.������Q1c���E�V�>�? Қ3{8�"�8����L�ݿ0�J� ����HF�D�}�A�"�L��,������bQx�NO5m��?��q��x��ho]�;������ ���`����i�f�GwK��O�uV����ڲ}^ъZ�>2��W��Hu�`j����?�������uU&u���u�cBB	v�	��s�^ɜ*��!�y��b����#�ü5��ޠ����W}49j�It>��$ޟ�4����	Go�\��t����~���P���0n�|�n�*����Qp�٭�Ƒ˺��=�1�&Y��{�	k-�X�����H�o�-�e���diHAD�9^�8;O��һ�W�3y��*Pc9��iN�&NN^��.�'쾉�Xp�r�yK�'�S�_�n�:L��P!��#�(%w4�)jf����҉����Lz�d%Έ�6KT����y��I��A�௓]��NF��?T�)���o��bwM�	eXc3D�v?kc��������	�xpQ�||�� k�4H��h���{���I��Pcr��C��tֶV��n�=�W.��8,H@O�;�z�#�F��'}��@�dM{֧O 8�ө}��GB��|��*5�iI�u�B+K�ЦW��T�֐��d��)�i@��u����ǽ{�%���XL��;V}���OuI4#|f�b���G�T�7<���`������+��#�N�x)�������1�B����".����Zy�6�/Ga8�؟�f���f
�-�E�0�o�<R�w��ɝ��u����C������S%BUmJ`ؼs�X/Ǹ�<�verw�9��-H�P�|Ҋ��M�/@�S�{|�(@~�I�m�QI�M���Hy2�¨n���ʠ���(����E����'�*$����c�"�G�tw����e6C�%v)�oޔqj=���>p3����hJ�B�T�qH�� �����w2QX0~B�ˋ���j(�LJ�&��xE�i1OE)�;XG�i��C�_�H���5���%7߅�|D&� �jʜ�s�V�s1.2��#�O��l��:Y��#)X�ۏ����^�l�7 ܵ�����	�ZKsL��("��+|�t���e7�=^������L��z>��<���&����+��Nzk.;�e�:�^=�^I�˩5� >��4(O��{5���7��{%r�<EP��U��3o3��~��+��h.+�r
"��e	5�|
��5*҉��O;�Y�,ߓ��z�o���|Vjd�����o_�пc�^��,O��75��"`n��gz[�N��Q.{�@Z�Ίԍ=,b2��2��9CD�m�s���ط�˙���Ͻ��{��뵡���O��"�j�?����|F���Z�]�Vj|G8}�C�?�y�~0�����urpȣ�<��=Gz�Ma�r��ɚ� �4.a��&�C�_e���e/󱐌�_��,*�ɷ��Fx�F�J6bP,`��c���Uu T�(�[)V ��e�^����&�9�Up���7
��&JJr�9���Mp;�=G����Uq�v��eR�e771��b����i��
[��W�߫�?��i�6<lh��"��߻���w��a����h�	M[a�� q`��L6�ɯ�T)�����$c��$�X��#�`rR	���n
���G��ϓ�{�j����������񝇊�o�k��~�tY�*�	t�h&/;;4;Oz	R�,J�Jk����*3]LM��[iC#��}�F���`�aќ�����l�-�;�r\�bY�mn���b�w�H�*�b��f���VE~�6�s��R3T����PA{q��䪤�.�6���ꋶ+��M*�A$�=� %��#T�r[1�>ة��A��������ڍW�%��b�Q5�ggζ��[GT��%���M���h��q	�]��;PZfX�b�J[G	aW�Ԗ�A���6K��u	T���^��K����HI��!9�Ւ	�2Ȱ8U�}��jzdԢ���*.��nu���:���b�Ǯ��s�H�sn���#A����1"��wG~�7[i�2��p�]\��q�����e��wQ�R"��<�.�Y7��i� &�Z=��cz�a�$�J�n��f4�jCb#�ʽ���J{<'?��ԙ�D��#��Cu@��
c���5�� 6L]}�
��ǹqQ���|Pp���O Z�d�z0�����Vv�dem�q�+�Z�v-)V'Q��\g!?}��L�Z�t���~ ֽ���y�H''÷�k>�,T
��B�Y�MIR�����x����gAzca �����h{ �k�mR�H�IL�>�>�03�NɃ@B$�Zr!u�|�oJ��ϲ�z���Z�O֪�ZQ���=������SW��EObi�0bin�DD���'�x�+~Xӻ���{�'	�M>��b��"�����r���o�.����� ����7�V-F��,l�1����}g�6i;/�!ˍ�B�7�#Q_Qђ9�Ŀ��bN�Q����P׽�^�vo5p^�� ����M�������@p�"�)�߮7�=UO��*/a,z#muRu�5ϝ>��?Sb���ls�<�W��g
�(!W>N�R������3�u$-l_�:�D�F�p|dļ�e�7 <��B`��C�7�և7�'�駝���c������N~�<n���T��)nv"*��q��`�p����1�� 
A�E�X�Fj�E/�;�X���>c�)�e�h�nfθ,�gH�-��@�UyVY��� �����z�njKݡ��� [����q�~M^^]�7��/�<�㒖��&����
X�A��
% �a�#"6Y�����|[����7r�gβ��V?��F���ǥ�5MG��/��7��%����'%���|�EE�����v�� ��x��S2�ps�O�&�n�����;Q+�ݪ����r�؂�z�\����)9�d�|�kd��[���o���M5�y��hZ(mU�{���"���Vod%����`t�E��'eH�J��v����G�h�E3y�$Z��i�N
b��n�.;��̟>���PU�k&�ل�	�+���c�}??�˗��?�t�1鍾"�mm�������;�P ������
ğ��j���(C�:����J	�0��$P�\��t����ԙXV�q��뫂l���t�̿�v�tm�<���u�ģ�/)�����l�C��d�s�؀Q�mhi	�,h[+"�}��ң='�[��-���u��#���K���dL����j|X����� o�
'�7ߑq�o���<���A��\�aaDS+Z��=n)W��������J�b���U]��fH������~Csj�_�Z�nɯ�̓�}�HFG��h�'�n��w�DZSg�̈́�I��3�s�D���D��Y�v_r-���ȍ_��@�F�xn|h2���f�)Ĕ�k���S�m�ҬFIR��2�Kj�	$�CL�Y,��M(Ɇ���q�Op>��QH$'%大�����������KH{�l�i�����dm���M�t����b�*�u`�o���(��N�L+�O��u�A9X�9�B�11�d�1ƞ�ᰬ�
9�� �B�0��қ����X�X9�������Ⴙ؏�ۻ��b#�&VVb'�8gS�Ft[�x̾a�H������Jg辱o3ԁZ�_��%^n���N 2��j0�}�G����Q��]�u�Ժ��X�?�?�>&iFAäG��[�B`*d�i�����DKγy	ʎ��.�2����(*�ԧ_��aa���%>��/٩�8}RL�HK$dBY�!Q�j�1�:o[G�X\o௬��k�{������_5[����xB�	���]�T�#uQ��7��
9Z����QRǲϒ!T�7��Q�&6�o@w���(�z_�����=�Y/k��U����h{&(�^�;qI)c��܀��_T�p*R���`�����3yu�BuW��CBy� �'�eO�>$$�1�:�]�C[��_^�t�~�6�O�*�rT�F����ńA���
���5̈��6�w���A�>��RD�(W'x����IxS�x�-J�HҾ��)C����)��닉�k{�T=&>7��`��N�)��O��9(�VW�>�>�O���7s�h��I�l-^D��=뉨�(�~:\_�z	2�����6`��oQ�>�����rH���tKȿċ+��&���ƍ>��=���[��S�W�@�7�et������wΊ�p���>a!�0 5Z~�޷�Y'�$��`J��K/�����}n�R��6.��q�<|гU&�d���� �f�Ρ�F	p&��j��e�*��t'�d��_[��嗻C��H��"̃3T�u;���i�M8�B,��:��ji@�qn��b-�bq4F�Gl�kD����&'5tR�й�?T����9P1���܎���	ed��V4(5�[8��U�s�t�&��Y5�������@3]���;��U�V��zw��@��!Q\Y���q�?��޹/(�
4�<Mn��:1��0�oϳ���Q؆�������M{�F	ѣ �����ɣ`[d��.�ڂ0�l	)��ި�s���ūu&������a���r�I$�q����'�h5~��&��¨.8>�Jc���a�'�oE2#j�����"#S�ܜ�4JW���y�a�j����2eU����1<.J�8q�]�~����YS������q3F��A(L'���:��Wb����kFt����=b~�#��C�%(VĻ���q��g�4^O!A��\(�}+�X� �c�m�-)�uY���l������t��g��9���'.S�b*����M2!��d�G=��x����)�[��� wj��=	T(sֆ��6�ͻ�2S��MS�~Kym�������5{|�hv�n����c��~el�kt���[���U2!JX����}�k\��B/�B;:�%fr����E����+E|��~}"��V89���yN�W�㢹q��p��i���Zf�O��J<㹤Iy�c ����t'/�7J�GQ������~�k�1���;�·�0�ww�JkIΉژ/��X�3��ߛi��F-͙!�>�����I�O�t�,"��i�2�?J&����y��.��_7
����Z��#*tǯ�n���d�+(.�>��W�ϱ�#��x����/x(5��e��N�L�؃Z�*��yTQF�^���+��d��c���t!?�؆!�����.��R��q3#c(�A�P}T���8�YÙ㭝}���u7�vw��X�OF֗D˯zRU]�J2�����	.�k�����7��d,܄��]B �7��q�4{<ݬ�X$>�9Ua�:�N�`N�K�Nx�_���&Į�f7nP.M��p���B����pJ��@���!M�� 	��9������d�h��`}p�xr�P�ռw����y��^�-D%q}����QRH�ӈ��z��C(�b�B/� �����p�r�=���g}f�M�{�9jp�R%'FW9h�@�DF>>��˽Pu������H���li��L�b3���*/�,=�{c'�ؽD-ë,"�cS]��^F�ֱ�|�+Ц��Ih2m�����y�����h���,�� �w^��(��r��B�fz�\�X��3�N�B^��dH�����!F��k��z�l�Ǆ��R�ﴌ��"��ja���U�_��}�Z0��͖0���Mc��˙^{o�j(��۵��А�GJ�6b��������*Q���E� &.��'u%���7���c؏�vv/�ɔ/�/�|�O��ws ��6갇x���՛�����d*�[��%�D�]u�]nnb�U���I���a���hz��D?���4�eܨ�YyɃ����OdˋriΪ ~��~�{��I�B4� �wE.�40�/����m���kܿ��S&Xw�F-��hKM�a<p��W"Ȧ^���"�}����1�ReT�B
�w��]h'>}������io�����"\�W���M��[�n�˅�l}��r�`�]��߹;�	,E��E�O<����\���Q�sC�ĺ"������_�l�fA�Un�qj��Uf��In�Q�� �U��WP0a��^�}<�p,s�V�	��QN�:��f1C�DV6̫W-����(+�,�������*��>s�W:ȉ���?\�I�� �j���NA�D��¼_���٨�-�TJ� 7w�L��jWey�Ue�D�g�d
~c�=M��8H�J`��o9����XF&Y�x�x'�he�㴾�;��"-��z����|R(}=JY�<O%�0�ׅ��m�V�� Z2Oy��^�ӸnZ����vQ�j���ǳ��=ߍ��p��?��r�t���ӝH��/::�7��6U�) �5�t0�fD4�p�{�N��h�P����Um���vV�0���}������])���5T��<.��XRL�wZ�l��^�ܻl�\<uu��hX�J@��aV&���9�ql���O�	\�:�vMM͚��@���䆸�t4xW��~5�{^��\Y�����X��l�LH�R�ꂡK�07_��$2��N�|��J��N�l0�t�Ib#��p�۵�o7��8Ml�y͟�b��z��VT�:�k!:q%��خr^��4q/�17�f����v�WB��#)&�ݡWj�/P|Ȫ�E�E�]��0���I������ʢ�0�_�h
<A����]�`�S��K!�V8uB?@^�����\Mڶy�m~^IHi��J
�����r�(�|fHt�5HR�,�	��Y'ʖ�$��ՓhS��9�ݹ�6��C�ψ��М�5���.��4#Z�L1��e�`�l5�r���C'��yB;�>׫�م*�s5~sH8N�b�W{�O(�ƿ��jD0����ݚ�c��׊e���t�k�������8��Q/�z��vRkk]�����7ߍ�/�&����Q�HY�x��J�g�Y
h���b��Y��s�5q_��7g� r��������(t5�|�@\/ �Y�o'�7e�s4h�'y�Fߛ��as]RXK����>o��B��k�"���2T�� ����/��t����P؎d��{IHx)�H��mYm�p��c���[ګ�sj���dnwP0�M���M
��<��¨�c���6�H���dm�Od�����kA.c�T�7o��x�p��E6N�Ş�)V�'x�E�p�����-����1l�a�t�.kS�ܦ���^�~�!��� d��L@�ߏm�c�R��^[�#����|�;֕�G˚Y�Ϗ��	�vP�GG��F�����O`���Ӕ�]�͓��NMO7����i-.�s��cǒ��^�@��{
!N����-)as��Ň� \ ���M�u����O0CF�)i�>_�Ul^ao�����Kl�*l�艤/�۶W����&�LT��O���n��Sx��YYw�{������7{�g�:\]��Qk�;L��=K!4�����5�[[����1�z�_��3K}S����Žá;��	�g��8Ǆ��_��/2�����ꨨ���CRJJ�")�-�(�݈t���3��"-!)� 9�    �� 9� C|g���~k}���z]�9{��y��y�~�9>�B�PE�/��~����B��z6=��[������YcAHZFPE+���m�3_���}/N��ɮ��G%FUY����͎Q̡��̈����GS
�7s�&Q�p�Є{�ڢ;p:�d�J����� ��U������>�V��ރ�eȢ����_fF`⧵����}�o�7&W�RF�s���8UJ"�e��yw�׳b�����i@�WL}�P�0���;��(2�8q"I�hR{��y��-t��P<m����BWUi���W$�����s_��-�}�<��jb�����Ź���\�h�OO
D�t���S�T���^S�W�eˁ��7jxnV�z�r������ؿ�m�k
%�=`�u@2���F~����aBʞ��7I�Nc���pP^�|F	����C�~���R[SWr|��3d�rN�.�J05�67w���R ��X����n���`����q���F���@�C��<�1Uk��?�|�ϓX1 ���M�7�=��k�\�o��>��r������M ��wk�0�����%��f=�pA_H#wO�p#����ވ�+k�(X�,O%%�p,��R_�c���׮vq�Q�Sc���*���x�x^��.�P%��41W�SE3���ƪ� �|V�|6�=��E&j$.����j�`a���z~�
��t��0l��))���x�Dk�T����k� M�ب�|{��<�	�%��J���&�~�H~u�{T�6�@F���u�c;Rgɮ�:i���Ղ���Ћ߼�pY��9o�o� ��Iɚn�UEg��Ǌ`�������f�����!I��T ��oë��bT0��b�Z�ݪ�}ӎ����s9�#klbB	w���d��y�'Qm�&)���/D훹�/���;*���k��w�0�����Վ\�.�k��.ڴ������ݥ*RB�<�@y�|`�����pa"�v��r��Y��������-X��I��z��m\�� �zgY9gJո#{�eE����*zi�G���:b����j�'!,i�p�K�8st)���.����H�-��E�� ?�9���r��x[ٺ���g>�l�k��t�u��O��l>�%|�W�j���lN�6�E�������i�i������K���c  ɞ��"�.�"{�Ȗ;�[���
����K8�/�����0ֶ��4j4<�M{;��)��# �Mb���~4�����`fe�nQZ�B�;�����:8�}^Q�[+b\.E��qN��k
��B����冣�\����-P��衽��r����B�:z.L�N����t���H�d���������#UN:>u����ą�=e]H����5�?7�p��Wa��`�r���R�Q�
;�x�L�SO��0BO��W�'�XXb��q~��#�~����`~Fێ�:m�.��T�*C�t
?��t6.�S��	���=��+#�q��F��`^�w��;�cj�s�;�`ȷj���֔��������oQ���o.椒��ZS���tL�9%u���_
�������<$�t&��)з ��yƯ�E��#7�j�0N#�sr�p��c�+����=*�Q��>��Rn�G���)�N��g�HY6S�Q��66lB��D�m�Kd&6)��'���YcaG\�~��A8�����9pu�5;��F.��j����w1�=L"��C���&cB��@��ZQ������-��$
"��y4��]�T`Y�����Zh��ځ�g�ô�LBɢ؄D��VY��r����y��w".�5x�1FUo�T|8�tLLrr|�zst`��1��SI��i���;��$^\^��� )R�C�%z��1U�&T&*�=�BW���6���k|T�l�Fn��
N�L�zg+��'�*ѝ���$<eB|�2�O����bK!�:Ĩ�WnOm=�����nɊ��5j�B~������v}ĈOt�vg�p�颫��iCa������0�3Ά���g	�џ��5~ĳ���7����t�"ID/M6��a$N�p�.��|��
Bl$���\1t$�L�!����	I�� b�{Z�>��ό�eX-�U��H���L����&8������	�<y����˅�S⻨����oڧ�t�� ����vt��#m}R���oB"�I�����{����JJc�ՁgV����|�O�%9m�q���8�k]f��Y"�
j>˰�ֲ�W$TV�*��^��)����I��b#��ސ�~�����Ol+���O���n~�L�74U���$�����ʫ���O�����|�*�[D��i�z��q�o�3���,c��#"O����/������vʖ+@�
bIket�������qZǙ���J��j8�j�-gF�Vl^(���ߗKJ)�t���]X؊�WJ, -��WѾwo�+��3s[lJL�z<>1n�1������gCw�tf�̆W�@����~I��t�_�nn��.辵� ���q�cĞ
�h�TQN��~�^4��x�}��S{�q��U����Q�U|ٱ��Wh��g}F�Zh�-����ܒv�Q��0�m|?�����g�Ʉ=9�͢��Nl���eˑ@�}����J;�~l�6qˋvdf� &4��J�+zä�S��ۻë��|���l��������u�$��%�����2����[����s��JDH�p�����Wǁ�ǧ�g2�)���% ����w�`*�5��j�*-����k����ӊ�?�lH��lU���ϐ����O�T�%����n}Ya�"a�#+�C�T�嫇�-`�،y��/�	g��X�1 "�,ʼPP����J����u�1�zd&u��]����95���Q�,�w��7/f��~'ݎ���b�a^���͒�.�>l^�n��Ȭ�fnO�E�z�A��2/<�	p���{EA蹌)Ɉ�c ɨ����O����k����/�*!�+XRĴ�'�NOFn�E=ÞbtC����ǘ���J�ts�5K�*�����CeR����XJEt(mgm��u}q�����Ug��
�;z�8N�9���{{Ka���>�ۺ��7|����d0D��HI�o�PM�N�M���]�L�o����Ѽ�nt�@{\I�'�Y�/�a��w�_E��Ȟ����_�B�5]�b���xf�h�;���Y��a���5ܴ�g��v5�'8���w�#��E-Y�	��WU�{��h�M���UQa��#5�F[����A�n�N���	F '����:����&�y��.\��0Hlr>�il^֮o�Wݒj��Lm�pf��n��A�U��d��שDad�2����Z�Jg��{ڣ���As0�;�zy�_���:�6���ɦ�5r|�B��#�<��$�m��&����K^�rYЌ�#�!y���f�Nɝ�tT�A\s�uּ�z	K����ȸ��ۉX�>�ӏLJ?�aS�P�j�&��^s�/��*�N��D6�w�v�]$��YŮ'G�����J�T^��)l�X�=2ʢ�u����*���VDm�	�{��gi���#+I�B���UE1���l�r�A���#w:['�ϼ�K�޾&��d������ϳ'������$��.{���/�}�9�C�S{�ZB�;g"�\�y��*����r1r�lC�@6��y�gX�����f�\)�q��ʹO�]%F�}|jW��1��ڒD�дZjY�`j���5����S�T}����ԀAU8�����?����΁3�=���w��W�j��sd)�7]��qT��b��HLJ�EE��}��I|�pÑ]'�b�_���.����PH�_�u{j׫"k}<��k8\})�'��U<p��������r�����(*��N�#�/�����th�*4n`���y	&,6��bVEa���$�u���w��N����ﯺT�2����w` a1"����������_ճ�,�=�t�1ޡr�=8��H�����t��Pj�N`�4�$��ǧү2�1�k���uS?cr�sw�ϫ�?�x��w��
"����~������z�Ycj��2/��)&2�'�
�'�L�Ʀ�����R�y��Z���3~��ձ��؈0�E[���8�֟���
����M��L�ݰ"s.�Ha�?̢�R/uNW�y�� ����Ͽd���t�n��6!�oRa�vR����\�Q�����9�n%�]w�Q�����M�Q�1m�
�1�-��5���ȿ�b�A���l_�F�ܵ���Q:u��n��o�Uc2�o�@Z�J�NB�����A�*��8���{8<�>��&�В�M��c��.?�B,g|߄�8,eN�}�X��X�?j������Ak~�o��a��"�X�{ ���`�������з���K_a�B��Rj�����f�yO$��; 
)VJy�C1�n��u���Rs� � ��ox���sb�u��E�b���ZC�O��N�{���22�)��,����(�~f��{Bʨ�M]6/Ɗ/�H쫐1��=�'K,��=���tv�q^���r�\, (�gIs�Ѩ�zF�eE���(B�ʖoV��P��HP��\w���-�r�6!�;8%���\Yg�g5:;���*��QD�$Dd ��@�,��l��[!����EIgf��ԝږMޝa,�0�/�в`V⊪ǽ��4�Yسb�z�+O�F��q���J�c�S.W�6���ΟL(�v��{ojwS�&m���F}{a���O�Ur$Ȟ�����E���1������%yr��1�����N�bN8�W^L$o�ǘT�����	�G�c�^Y��!!H3�Ca� �qz�|�W��o�+�;�U�:���w� l����͠{�����
 q�N{�q:����t�k��cf
"D依Ea��VU��z�	\ȑ�h1��1�ۻ�pnCja�_1�囱gO�G�L�<T���0q2�+�/9�V���$�$3�χ[]�7/y_�:F�FF�c�}d!/���z��r3}��vGg��z�ZA;r�Ǻ����[W�K5+^��zPT;鸬k��0������j��Y��l�c||�ar�:a�r����� VW���zaj��U2�̱
�=��|Ӭȼ�hb"�@�^�Fm�0��"��!��QR�bE�Mof�� ��l�5orB�W���6����I;�G�����zДx��
�{p�M���Xr��
�"u1C�]|Z��|9A�2�v���`�)1�-P.���	g�%K����g:X�ь�>,TU-˔������M�4[̭*�*,@2����ah�U�qؕc���ی�7&z�KiK��M<��8ڞE�t�=5H�E�|��d�0��y�-�W��s��{�6!�|��ˣ��� �p$����1 f�✦ �@J���J�����;*w�t�0T�=�wB�_�wڤ�I��7�R�z|>���� ǹ/���|�}�E�'t&5���l׏�������^^�x͇u�+l��U�y811��}�r
=��1���w�t-0TG<�7�9Ѓ���ic�`���>���S��`ⱖ$���u�Ԫ�0�xo��M��M*����^p�KH��;���{�L?�*���&q���h_)�V@�bǏ�2e�۸lc��K�Լk�[>[�>;m����9i0�r<j�K{U�6ѻ���bγ5�5�G�l5���ܤ��$� ��vh]��d��/��둪�� ��RXׇ읈��.��s�7�[��?��
M�ȍ���g��Aw�u�#�4�~g��Tk����>E�Ct�g�8G;�����c��x);�ɘ�������x��xV2Q�9�$u>(:��
��U� Y�NT�t~�r���F����@����H�@�^�_:���n9�;����L������ڈ�_��4�!o���KQ��|��しoUf!o�S����ӺeG�n����ӯH���t�����R;��QD�}��|��ba����/��#amȧ~�6�f���ӓq1ku��M��/�<MJ���:�.�Z��\s���͉��e�bַ���v�����H�g��n��ϲ��υk3J��#��`?������pw��.{XeTe1�zz�R��̢�@P�Jg��z�իN�\�b2Z��,�8�1_l�^�ϛ���wRBe�d�%��ѷRR�L���Ժ~�čǘ��x��kG��Q
�����+� ���8ʐ?/�M=)g���,<��@�Y��B��������r���ݶ�B&�Ю��WY��5ϳ�k�@-Կ�� r�N��bd�UN�Օ�c9e��>�U�S�M�G*�I�Ŏ����P/��k�䰟~8'$�:1��wRΫ���\\|���#�NkLo��������?;Sܬ�I)\ّ��Y����n��%����}�庡`
Z����S/��Qi��F_�z!�-�<�A˴wI�����s�S������l�6j�s����>��p&&
J3�W:M�$u�2�k-�cn�bO` �,���Sz�3�;�W-_�\�'6�i� ���x�s�F#�1�e3��:���y�s\1&M�`�Z�w|�n���m|{��ԗ�����P1O��N3��3�GR�Ľ���@�����1����ˏ���� <��AI�\m���b�}�K.�b�T�S��g���(;b�~~��>�;�����F��߶�����ep�MH����<j�l+5EI��{w�i�A�e���Qz���,�|(2_�0q��ycڌ'E[���+�U������{~��V_�u~L��(�]�+�����w�d����%���q'm��`�+^!q\���Գ�+��%*� ��Ə��/�N�Ο��i�=@gG9Gu� ��p]�5(�Z��Uߟ��©��é9�M��&i��g��3Ry/��w�f�v���[u�������A
����>	�]��+��g�|t#G�Tk�2�p��NQ5�_{��r8�H���=eװ��NՁ�23��q
�J���K�/�\=T[�!���T���tA��S6�bK$gr������J�y�b��F��k]�gj�
�o�d�#��HCcq�>��U��Ԑ�M��	
�������x��-m�|���^���kz�A�k�t��d���b
Bk��*������g���2~L%L��\����j����$�����H��!A�T�m�ϡ\[�z$L��J���\Tz�:Rc�����LƳ�+�lK�J ���3z�R(�>�,i�+\�SF��o�yD�\���=IZ�M)A�"V4�`~d�e=�Q�ŗ).�%������T_��Z�~�Z��d��"2�J��N�L�ю(��k����S� rașTy��R��z�l����Y*2AJd���tZ�(<[䓰G�i%�����N�N3�-p������]�@fD��l�ʣO|��v���� ܇����v�d��6����� �k��)���"��ba	�3�gr�Qҥ���1+���7�'�1z"YT$˾^
�ޗ�C��ֈ�77�%n;'���LHX�0�5����փ�#\��?2F��Ea�`�E<EE��8'���g�t���������|j�UCra�6�kNV���.S;/�#��'�������:���;�L����s�^h�b��ՕX���G����eϳ++�]Q�A��4@��	�:�ʟ)o���|H"�>m��A�I���,�^˖�[/���j8
�T"���/�|�$��͹��2ڏ�Y��Z?�;e��Qg��4�nT0�_%���w� Ỹ��u�Nc�%�^�r&Ϲ���i�|+�n^�G�)�&��b6�gԌ���Կ�7������9X~Ƌ�1�3ry�Mm��m��K��8O.�#�;n�4�tȇ]�:3.Nmߞ+x���� x�<��v&<�:����v�z�߁ؖk	��9�^]7�l�J\O;m��3�t7�;���vw�4�ţw�g[��7p�+���^�
<Co7ST�lix���$0Ya�(�F��X�D,<�S_��Uf�vA��i�B3�Po��H�/Z�����ŕ��-w��	,`��ԋ�J>.yfO3O�Y;y�zI��[0}گ�GU���^�80i*��[>*�/���+\� ����1P�l���ӥ������i��p���"ے6�П.����L�5]�t�� �6�<$n�)m�/c��)���G_���X�ߏ�w�:�=�m�d�'�.���������着D"��)h�<"�%���N��hh�Kq\.�ё��o�(�Z����䋞��mww�I�p��xֿw$`b'ӛ�6�o����4��t�Cb_5�j�F���N8A%=�h_p���5��-[V!��-Al3�ٍ+)��߆�gk�Qawvs�Bg~��'m��Mt������}�>�1�[0Zb@:00޸��p��d��ϲe� ������k?a9S��/��e&�����.>�)"�B�h{U�`e���k ��V��kk!��-�� M�Љ�cr �>%�z���o��j�����u��,��x��ͥ
�4J���n}v�v6/�ʎOw��,�u&� ��T�rd�;�	1�-������>��o$(��y�Vڨ@ޓϲ?����F��w\	r�{ LgMv0^��o5@ެ�\�����!*R��9�g�	��?LM	_3#�ƑKǧ#b�mz��y��ʀb�o�p�	=*�@����5/�c���ۓͥlS�	3�K.�7XS�ү�9���tTAhu,��lNԟR������n�;=Z���ÿ����R?��۫D�@�?bm� 966bB���aP���)E��_�!��f?[�X��{�S��e�u=7kB\��*�H�_%6�M����0���eS*�C@4�J�R����Q��B�1�9a��x ��i�
�ߡ�} MQ65E ���h��/��a��;����{�^"����΋�/㍅s��e9$	A�&�AM�UU����-|*<ch/��T~��K-����BoPT;D3'��O/vbq!��F�����M�BN/��Oo�O5��BG39v^Z<���������{<0��Lb �S���D�2��4NP�R��F�!$�j6%���R����<D�a����)5�Haӧ���?pvsT�M1�ФF=1U��B�5����ݣ����3(��HU��p
S�l�(�;o㎫�|�-�N��(��.����smT�NN����YK$[H�o>�m$��4A�C@+$��r��ﷀ80��44t$�wS&�����M7���Sl͔�k@��'�[�*O��0����6�G$D}�B���Ћ�^�����Ɲp�D�����4��$2z�W&��ZK����iX�G2<����%�!��m��@f�4����Ab�q?��6^��ז6 W��Hm�d�B�}�W{,�U�  W
�)�ץ��F���	�)H����C���DN�)���g~�
�n�r������K�zğ{V(�E�J+��[S$�;>�2ܤV�!��|�n�ǯu�20`��йR%�7O�J�<��vT������iEʷ[����gk�{
��<�{~�Ϯ�;�n���_]}��ߝ`L�W!ߧ����x� �L��yT��x�����w��n`�d]�U�r.���)k�tv��n��c�2ڏV� ��?�"5�6��:hŵ���q!��ԛQpp��
��[c�V9��G��cO���ߏ�ʎ0��[�ޫ�c}R�ȫ��Y_� F ���Ϫ���NA^�Թ��`�BtXA^�B�h����B��%����y�J�=��)쒱�r��"�[�9��1xt�r�wJ<�й��h�:���iW�p�9���YU�A����t��ªc�����?����p�Y�w���S�e��i��t���3�>�q��f�-8/q�����S�zl�.��"7�jEF��K��#��+��}�>ݜ9��t�6R�J�ݷ{�����Rqg�'w���@K�{.�@h��sr^�`aBf�&N~+(�[����P�����c�\��{12�H
��@�j7�������i_RO�)�̆y�=
��)��Y`��[{sO�(�O�X�%#F�6��آڟ.C@B��
��cMZ
��#3s|P���	8M���VXOʐ��^�;\�Ь�$�8�ͷ�"uʮh���z�>5�/��ه\~�e~_�q_����z���?��<PDۈ-��EvR'���\8}@���,n�_X���ߪ7`���m��v��/���n�ߴ�d)u�_�EU_D�����Y=��ˑ�X�c�u�}s��H�t<72�p��V�X�u���p9����9hu���� �M&�p|iȝ)o���`�Zտ�DR��`��Z8́v	�mkj+=r�q0�Y�<P��h��Ňp�m	��d,Q'�[SΈ�s�"��}I�����%�d����D��S�>�.F!ї�����'�\���@��p�̥�&A�GV�kkA�Ʒ�o����&$�I�H5^oo�ET��K4��q�7�nKmѓ-�n�p��8X9�k6��yi��h7w��?�i�ЙKy���Kr	��[Q�-��m�_�B��Fz}#������� ۫���A������ܕ��>�_RJhb�iȏ������VP{6J�+0/�__�O��f��Y������&���"��cw��I�>o��HШ�ۋ���Eɕ��H�j)��6*哤&ѵ�`/��1���):�y�yW�p9�����e6�z��GM��y��S�ͨ���,J�(7���[���ۿ�-�iͺ��V�BrU�G�VΝz ʴ�w+y�CZ}ՏQ�W��+��O�ߌ����CPQ1���D�3�aX�ۤΌ�Y���زd;ܠ$�(%
�92&n�e �OHv�tNT����r��h͐�ԓ��x�`_��P�Ḕ�1����*����` A�)>[z�#�g�#c	��^-+Z jd�,�� j5���L�H=A��]�'k@l[���a� roW�����н���i4"��Ƽ�g0.�w�&r��) �E#%��69o2��u�画0��-H4!}Ɯ[��L`��/���[p�ap�,�L�lX��b8#c����ZV�I��x��Q��Ol��Hl-�%$�_`�}���ܬ�X�y������硔ܾ��~W���c����'5��ӭXV��}���$�^��~��>�-$�=I�2.�Oy�^$ KE:OF��'ٵc �5��2�@܉ޏ�Ы�fm;�����T�mH$u�S�y�ү�S�|�Q!|-^�`Cb@.�O�~օQ�΅��\n�ն�!��� ~ H�����G_Z�/�,�^��M�3���#�g:S�WЋ�#�#gp���1)2��������`�Y�L!�����;��ͮv�ՙѮ��4���!�cD��Cy�h��/�E�a�L��b 9H�c!��=���n���e�юq��l)��5���������􏩃Ǻ���b3�@_���?i�������Z�xR�����R�w�>�c"���(�U.��푒&��.ZA�1qD��;
h-8�V�$�6!;�f��O[-�<-:�ͫ��\�g�ƒ�a�<]7	&X:����^<��{����{tBfq�eM0Ú땄f&*�TW�u�?� ��R��8�F���mL[�67t=�n��cN�����D����� �-yQ"8w+�y ��H7��^GN/�@&��emS�	r���J��mU��x�o������ ��o�s�W���	���qaP�c�� -Fn2��ꍚR;����ށޔ<j�W�4OL�HLZ
�������b�j�b�ni~ΰ�3���2�\l��l���[�J���۪C����H];�;��  ���AWװvWڗ����%�]|�3�����^�][T�v��7���_j�Q'�g.�3p����9��v ��;5��'����oIo���ؔ@�14��ǿ;B��i-O��ׯ����X���3��z�Й����]��p������$��3�^�{"|����j�[i�3?g��;���o*��"�م����U%%R������6�nc`x����IÌH�ו﷈wHpo%�O�@��Ҕ�� D�;V�.d�C�%��� ���dŗ���Q���f��7�<�6���ʣ��-�5��]P�jgD�K(�7�r*ͥ���z�}��zc�׌�����R����p�x�!AD�=���Y��r�Z�ٶ� ��г���"�32ğ���Y�j����)#� ����'��ک�#�G�x���~�!��]Q>�7L���̣J�`����:*�'��OM���-��çV�.8�#Y�Kϟ��[��_'m0�V&`���?j�,����ro�f3t�]��?dz�o�aO���Y�V±r��h�	�;�1p9�֜��%��&�()�e��?����.��j�+�"D����X���P�8|A�0%娆 ��#c5��%W�v�%���&gZ�+�H�q�� �e�[5��%I!������P>2gĜ-d6��1��C�;K�JsK4:��Oho_x�m����q��afv�#X�O�ٟ��m���U��)�I����Q�/��`o^e��y����5�\�������; �������P�E���Ku�ׂ�nхsa�t����0�ސJ>5f���.n�N�֐$ :��셈�*\��x���L8�Z`Ϛׇ��9��2ľ[{��<܇��2��07�:%��T��Y�G�fR��.��ES\���B�Qh툉��EI�痧���»���m!r0���R��iu�ϛ��q�@7�pd�q�ФQ@`&�j
!|��*j������Ǯ�����u�V����r̲<<��Hۚ8�O`��{t�#�85��/��ǉ�8��A����=_���1/׳pj�:O�� |s��o�d�.�^���77��&+Z���SJ�ƴ���J���N�W�R��z����''�O�X��P'A���n�۩�Z7��<^a��I���lU�����k:���*��Ȟ����P��=����Nj��GZ�A��cՀH8�=ݍ�QBb�Ao��L��cp�X��EY�.��=Ø�g>��O8���L��l�`�	���${BW�����Kw}D�kZ��<+]�Nυ���;]!["�Ϡ��B@��:�|聘xE���+)NA�r(�s�=58��1-[!�Ng���1 H�'��|)�M�����?�b����YSN�����1�vEx�sP.��sPZ��x������ssm�l����`������xr�o-8�<l�ɦ�}{W��LX�X�l,(9突:�o�6����#��kF�R�����q��"�r��2��	�h)!5�!�" Of�&y�� ���\���V����kd^z��h������A�OK&�B�x�k�A�%)���C�N:[���A�1}H)MG���z��X#K(<o�c�����ж������0qՉB�?�[^����@rYT��Gc)u�-3_η[%�F$=�����s7߹��զ�]��n���q�:�u��E&X��|ď�k��*��B��>8#[ջ�1&$$�;6�"�.a	���
2���kO��ft"��fe�~4MS�S{9j��;�����bn�J�M`9����r�}��#�+i.]�����>��KJ%4�ZJ�?C�1���QT��@��>�l3�~��!XO�o`
r���������Q������|d�2�x�����(�6��V��n?���
y9�F��"g����΁-x�q'�B�}��烳��C��HA�������F�z VAΥ[�4�#)�����at��@YT���������c����f�G��vD�b�����xI�`�[�4�i|��x�{�;����U������kC�Ho��FNj�������6@*�"y\��U�;��4��Z����i�g�N�oJ4	H5�"m�,MG/��^����^����v8��~4�s�tL\^ϔE@O=./p ��67����=���p!Gߞ�ҹ�z�N��Np�i�R�5��)�5���#�fC����uǅ4��ʈ;y��]��s�0\�n�܅Dbp�u
a����Op�9c�P�����@����p���⁹�K�Ƭ'NꍷF�����V��,i���X��`\��rj�;3�W]vU��*? ^=�����T�����F"�ޒv�z_����DrX?�>V�����5o���~�&p�����Aߺ�'R��p�"gL��gB�.o(��_i�<bM���F���B����]�]Ӯ���o�X1᫸�LD�V�+������R�__�wq�U]�I�2BB)+�{R�<�Μ��]�x]�H�nBm]�����{�ɮr�h����X��H��ľgƀ��<��,Ϛ���R!��+X��Y�d�9|eG���s�K>!ê��8
N�k��-�� Ζ�󭬞�����Q��1g	.�R�l�*��Z�U»��� ��a�&Xv_Y
���|��&Vĩ0O�Bg��Gf����GD�像�Boj8��8単4�J�͋��L��)����3�=��,Kd���=����_�m�Ʉ������H�_�"��:�p�y������c��{Gk:tՊ_ޞ�"�#��)����M�{V~HZ��׋X�Az,Hl��1c�߱���If�G�3C�t.Ժ�U$�7���͖(��ԈI���8��$��8f��ԗ��_�(��|~����e�OG�Eo$�e�A�̼�hs�&0f��pF\\k gq��t+	��J������0+wA��@�]��h�s/F��0a�8�2�R�-j�e�X����x�ѽ�	TnՐ��z��D���w.��rR��L-����@�ĳA�͆����o��]E�Y)��1��".�t%���c��4�b��0����4��8��"�rpvt$��'%��`������_�:��#�J��V.�nY�������N�q�?��L�7�P-I�`B`�N�:~l�,�F伡.����#�͠ �Ws�|``5幰�])��f��Ø���t�&u`�4S ���U�����}6�7��Ō����*�G���Ƿ�rᓭ)~V�'3 �"�F�0����Չ���@
70���~ȞJZ���j�${f/2V�xﲨX��j~d~��_�5ԭ��΃�@�;�^�#��|��bs����/�����B_r����;.h��v�����7�\��T�$Y��I�Ĳk�[����D;����2�N��ͳ� �u�՘gAg?R��t�̲?�/H����_}-�U郎�\���S���*��.�w�K�հ��쨣�ѷY� ���Nɱ��4}�b���~i-/�d�^�Qͣ�(uv��39E� �����5�6`�y�\���P���+�i����??	'�IP�M�����涚�eּ��,P��ޫ���?c����;�T������z�v� ����D�pך���x˙sy����mb��O�<��i��>j�	&�y�^�N�بgk���$�t��7r��J���\��\�յ��KK�
M�{33MPT�<>^���@�ۯp� ����%�vf[�)偝Ebb��o�ž�Vb��̏��W�\}�B&�'+�Bx�a���Ow�Ծ��o,�������M����G4���
ڝ�������_0G�����"��<�Q�w}g�Py��?�ž�h�sM�z� )\��<!l��B�װl>�z��PJ;\*r�ߋRk:?�����3��	Zm
{�7�1?����̱ٙ�ة�LtM��[?I�/h�W�jI���@�u�;�5Ew�z
�^�� ��S.}%M�6�)9�w��}��$����o΍F���LW�� �L�zń^z���P�q�⺵ԕ�+H�Ry���@�[>��Gv�L[�(�g��;q����?R�G
X�-zE!^>�K�������{�k�q����%e�1�4�Q��h�k�;��A�:�pb��l�8�8dH+UM�O{���8(��sb�G;b�N]�o�l���>�?]�[���]�I�(��Em ��i��G�\���uc#����U�F}�����b�i�Q�>	H҈ɅA����
*�O.<|�f����������8WZ����2s�^��ptzt��xؒ��/'cY��z�$���x��\�����嶐�G=u�A��)�����A���oȵ��5����]�7�
�.a!��X�N�I�{��t?�K�;;x�hg7}��2ᐺǸ��ׯ&�]�oG�Q7�v]�ŴG�%�U�i�{Vjp������xD��u�ErvR�Y�� `?AHid�,�� R�~�I]5� wEu)����^�u^I��V���RHFM��r�R_j_�-jyOW��U�k��W��+��5�=���X�l@����ۏ�1�J�C�o������a��l��d���l`�B�{-V+;�
��L��5��C�3愴����Q�W" L5EŽݘ��U��w�/�%�4_Y1��s%7ކ�R���0�I��^V�L�Cu{*�v� �g�+��w����3� !�� �c�n�r��
e�ـ]m��m�Kx�ir��Ŀ����%��`�#�@,�G�!��tEvYd�p'_2yh8�q�q�����HA�P�����tF]@zgΦ���g��&,��ס������2�i�t�L������mt���x��$n"CsO�e��!x��CWdU���C�Ψu+���u��%.��8�7m�i�4ҿ�g��<�)����l�o$�����K��a ]�����P��t�X��2��q���*S+��]���m7����S�&�'��8^��Q/��x�1<,S<�>T�5�^>�&J�k|̻�ru2����m<�2{�ǃ����mR�-���Gq�{ܼ�������z�޽�%4=[�[98�h��W4�����'����f���U�.O�%�6�4�56tL�}�n%� �̶����m�%2��筰3�uX=�$����k��iJ��H��ۏ����V�z������:�3)y���$^9��g�x���Q �3�;�3�#F��΍�f�4^�;5G��;k9%&�> y�#�h\����B��W�}N=tx��
ĩ�Dj���
qa��&���D�����aM�]�p\��Ea]�""J�^�G���ґ�Kh��(u�5�D@@@zOP�K�:��BK��L�}�x��}?���t23gN��}��Mfr��2�Tl��zΉ}^�S�j6�u2alr�2�X˕#��������L���'�t�@�n�ʀ���iq���@>Z9N@�3���6��h?'�Ӯ&a��H�O	����a|gO��\E����ʇ�q8X�9���*�R������ӐC�1ev�)����4�X�o�9�K	���!
+�WoO�l~"|:?p�s��Y�ȫJ�{�4��yz2+��^WA�
eQg���K�wE�V�Q7����sH�._-'��/ �^\�5�󹾯r��v�yN�>{��M����Ҍ1?Y��X��"2}[�~�ҭ=��t��f�D`a���՜��l.��-s\QY$�KJF�٢�ܲ7j�Y�����8���*��]��zz�.�yM����=����tqV�����v-���x�{6Z��ʗ�̝V}�A:�OfV��>yf�c��5Bz]jm:��ܹ��|k�Z㽫�n�� $>}"u����m�����pFf&�;6p�����Ȍ�{%�2�&8��!���a>������R�c�Jv6Jv�dg��Hֵ��d����3[U�`(�gȔ�����������fz�� Y�E���N<CS����=0���s��~���q��ʵ��Y?\i�u�w�*�8`溯8��`�K�M��ޭqT��᪡/�u&]l_A�X���e|Y_=i2Ns��i�������Hc<�n�t]��K�Z�3��9�;6��ǳ�'>��:χ�,+��ȶ0�~"2�8��:.��R-�2�Z�#��|��ҋ���+�o��6��l�>/�Ђ�w��,��}�A�@�!�xb���c0+$��:�8�Y���~����1�=-�V	���w����%u Yx{M<�2�j%W}�{:�1���d9��$ĕ�X#��²��:+��I���B�</8��Ռ����ȸ���y� r�O1��d��؜�L���fzg�~W��,݁>&�~z���#^�5G֐�[���#6{7]^N� ���w�Vp3�X��Tr�Oʫ����z�Z#95kē
0�镃�	?�78P�==��W��3us7�I�ە�Z��?qM�"_��H�O�e{�0f�t�bf�`f�����pn�����/E��?�e��z�I�f���wŗ�@:��N�r�H#�2�TJG�|X��R�O��!��@l�h8`�BL��e�vC��Yi�/޺y*n��)t-��₨G@�1�1r�������~�ͣ�1��n[��Vz��T&7 M�o�2fr2f��4O?��҃<��*k�j�D�Ʒ�_)�?�E����B�?m����z�x�TNn��i�N+p��%��m��X�>��B��`oq��T��l��F�nL�6��N�ʗ{�Én���_WۡBPg�����6i堾e�s��#e�Yj������E|�*m���4G��ϫ-��;�$�;p¯[����ٗT%���c�%��P"�"cNwbp��K�����(���E=��]8O\�������������嶟��K��b���.�7�����n�j޽k��Ok����������S��oz��jߛ6x��X@?���t��E9b�3��Ҏ�������S����� 4�}�]�7��B��A��6+�&�О�[��] 4��；��c�T���ESx�
��
{����Ș�Y�l�3�Uos���w:�^@";S�k�q�쾮@�X^dK�OAt�����]7�(Μ:����C
B��ʧM���)�a�����Y� ��
b�5�j�8�	�	�SW��C���� ��Z��^�b���•�L˽��S�N��'/ĝ8s{j�	�25z�O� ��3VR�������G���@J��:ޯ/g0Z�'�4��*܍)�`�EY�`��?3��-'�k7N�66�)�z�uQqϯ��"���2���ϳ.�}�d��e**EV��	� ��t* C�W�$a7R_<�#!Z��w��l\]I�g�	a����o�@J�X�vXLt��R~����n-k�_?w��K5X�_����c��>dx!�R/�qt���%��ޢ9crc��r��������ڧ�/Zj��|��"U�g����"�m�%Wֶ?�nw���x�v_��.@T��J�?�ܟC��:����3�ţ�|�Ej�F��#d[�孏�|N1���,�v���gw�l��!�<ǀA�[�=�9m3��Q;ϙ�G�f���u���A�|m���;=wý����3`�5��`#�qO6���_r7��}()��cOm'��NO|���?���U�滥fvZ��%�1���� �Al@�  J�����t�5o��V� �˕6p:���Ѽ���!��O!V]�jN9m�� 4m5S�FE���J�/�*���̖����n?���Q.��kk̛�~ԝ�H�Z�����b_N2�^엻�"#)Ȟ��p�˷��F��>�x��	�ష����u���R�(6O?��7��+�����L��Ypv��*/gcO�O�kU'�UY�����U���2ڂG�����K
�S�b��r ~��Y��u\l�~A(5]�퐡�[]n}Z�qʒ?��
i��`RN������_��i���,��yO��.�����=Y'��9ؕ53�n+sU�^�;��p2(���Ĺ��8�q�sF@����'W�d7;�#dw;U�r��i�Ͻ�erxa>$���9@���yOy>���ߡ�݆S��h^�hx@U����dV�R��H僘V}�t���ⱖ�8Ks���E^��Ԕ,r�7�0���|�W����2��F�������|8o��*��덻"�F���I�Ĺ�P�l�,/��:��S܈z	�̒t�×���\����9�d�5z����Լ;�q3��sť ۵�����8���ŝe��D6,�������|�Pw[��T��o56���khRGr�H4�m>`nJ��G)��`����:�M�;М/lʏ(�RQʻv�@{}�4Gs�9P菇�2:�I�ͨl	㙯G(��4����z��J�j��7X��{h(gF�[C?��8���������Y���![a�%sU�Y*���ʷZvf�oL�c���m����%6]��Ļ�d_ҟ1A����l�x��
'�p��V�KŴI҂#�-�u=���'��f��R�͜�]��6�2��.�;���w��
hFH���5�2����g<}���~x��#v��t[�K���~gR~�U�}/��/>+�}W�4�Y�u�y���5��*�@?�3��P�ZcՙW�`� v#@dn٦����ZԢ���.2�:yq4D�c���2Ax����Q��7P�ag=�Χyu~.�7�a�Q��Ө�]x{S��M�۩� 1�q�+ot?�Y��c��t'-�#������k�]S��
�ͶȬ�N��Mv��s��t�n��R��p<\@^\P��
��������a��������Vk�&��ai�]�H�5���[�f����L�$�� �xb��;���B6? C�r���L�~�hG
�"PZ�<���fo�Q��2�c8�2��D�)��X�����=I��vo^����S(K�[Ăm;09�M�Tr�<*�*�T{�� �|f���&��j^_w�|HY�c�j��Z�l"$t�D���j|@��~� ���'=��r4�b�.A�!��#x��1縦�\3.�#�R"]�����?(g`F�l�w�k��+e�c���olb2�B2	��"�שB��g���B�����$�Yce��|@������,)�\��G�w�zw�X�T��8����'¾8�H�}ac��o���cL^�)��F���|檝Y��r��G�V���ņ�[W-W]kO�.u��:y|<K-7���ty�Tw����`ݟV'ơ2<v=�w��PX��������(�^��q�ޚ�Y�����lRl>s:����Hb�g]3�bsn ��p#��f\zO�N�O�eo�0SH����;H.� �z �ƎeS�E1s"��2�~��e,qi���̞7z�����9/�����W���<,b��4g�	���R��Y7������3~�ц�h?Z�%��b|�m���$�� �����B�d���Dws��ak)�p[1�Mz|�J�Xi��=F\Z��^�.�!.͇��(��gԷ7������̾+8/^�k�q�(����]�U�TZ�S�l���PK����mȼ�$h�'�g����=�`��q*^����N��d����	}�;!���A�U�8ǘ6ǰ�:SY�W�=cf�{�]8i����@ePl*&ȇ��n`�J.vC
2�m0��(�hbcc;����2�?v�%J�i�'Ԏ����Vz��x�3VVl��f��Jn;�[��w�5BQQ���Ѹ�:�t,�~Oz��}
��͘����̀}�sY@�4�Q���$ �ݣ���-�!�1��i�J0bR�^�Ɩu�!u� ��=,s yI��49�"(Ή�ZtU�뫦��"�k�������� İ�A�W���D��_���mݜ0�z�{�9�G���� ������j��gj2�����l�j(�۵��� �P����̹[�܇F[W�.ܻ
��{-]�� .��MO&2D>�5��Z_-��>ӂ�vE���	/��|��"堬�Ƈ�v3��F)E��Q�L���F� dkvr��1A_�) �������'����X��@��p��'Ov���;/�1At=�-U,tk�� p��+��.l���`�"�2Z2֥�h��$�Ǿ%�����=���=�~y�?�̙��������%Ģ��@S���ӛ���>�J̚Ԛ�{f :Y������+�DiP���W���?���AAt���̲��4�C~��C�"�湛���ư����[͉�3�t�_-����ô��~��H�_�$��l�h���20K�A�&n nV%S�{��}6�t����SPTf��<���Z��I����@t�G�H�y��DC�GȬq�jď8���*t��D3�/gfg�i%�n�,��ک�w3G%�n���|([�f���^��9K6�[)����&�F!���\�N���V~x]cq%"3� �ڦ+�H�Ո�x�:#w���B��E,�,PW`��R�����^�᭍�l�X`��S[��'0>=�����f�I�����RĆ���u_Azgٞ��$����{i�[s�7{��17?�|��"����wF�!�������8���
M�W����:So�7Dǫ_�M�&<���eC�˳��lp���X��S~������Ia
�404��|7�1�KXR��TDD����0&�"��(/�X�qQ�Wm��u�!�0�;��
�2	�h8�\�� �lm��0�ww�S08�1XL=�a}U�;�S�뇭��9+���K��+��F^�����˗�{=�:�Lj�
����oЎ��N��z�����$ō�j�;�Vi\�qJdF��"�[����
�� {���EԚ|�[�ž[�	Ӿ.�G��n��KKp��,	~% t]�Ҹ}9i��L��b$��b���m�2|�@fв�v���5ZfJ�}����T�X���u���B.�fl��5�c�3�=\êӃ$!�Ǽ:
�;��T2z�W�~��RZ���{Q���C+��HhUV�jʲ�݄h�s��׋L��W���bh}FC�V2]�I��&�؋�nĨ�o�qpP�Ɋv��%��b��P�mu��Oܙp)�IrKr��SFG�q�[>���t��������0 ��9�����e�J��[�4^�\��0�c.�Q)�hoʥ�?661t����
"���4W���?��3�z�Cxnжp��܍��Q-��_u]����4s��w���10�v��՝<����@y�e�#LW�QgΪ�u����z�J5 )�g�޹���g�*S���I>�Q�N��C_z�3t�5��8}�|f��ጧTVM��=H� [�R�\w�g��_���Bޔ���G=_ג8�E�RZ�@0~�W���&�����~��d�I"<�su��_(sų�Ӿ��w��K��`�b�H$[�N�l*T��f9�͚=K{����
:ss�5�|��8K�r9#:�Z�����y_H�H���Տ��z��6�W��QJ��/`�Aν3F�B6/��� Wj��u�'��t��
���� r�S��MB�+�J������MJ�R��d� ؓȸ�\;{V-B$L�ӳW;?�EQ1s����	~�<Qq2�lrs�����3��3�[���q�,
(�����2Kog�����e�-�ǹ���k������u����;`�ǻ[�(5�c
���D�C���]ͣ$&��
k�8�v��3�u�ϰZ;h_������t{��W��	��H��Sb��q�ga0z?^��A�s8�w�03�ڎ2���ہ1�T�*���*kP��P�
�z�48��.ј���t��*aO��[��H��-�9X4����;aЭ���,�:*�,����T�>��bY�У�GYl�����&�%�ǰ����{c��XU�ږv�9;�9���ip!.�')�֛��s]c7����8g�QU��{7㙆.i�
4q.�P�4JBWV��| S��l����Ϥ�`\��M&�n���i��%MW�7�������>�3{#<��\]�c��M�@�/z}�OҢeg��A�1z�,6�57�V?��C����q�?6��6L�+��N�'VGA�oWj!��Z*HP��S	�$b�2��o|��s�DV=f�9 wBe���8� ��ۜ�í�4&%���~������y���#�>@qډ��Πǲ@XfU�u�ស����YOAR�'å.�11�>��L���0��H�q��U�C'h/���AN��OSO��������dxM����(!�q�I3���2�F����}��=54�[y���{�j�z��C(T���B��~����w��Wed�Ӫ���e"(YA
r�U�]@���xV����6�E��i݂�P���P��B�"�@��Gg`���� .hR��� �a��{�n�|�߂�z�ޑ����◲�;��l]0�=�T(8O���$�u|��J�� .�B��,�[����W*�
�}/ۘVPQ�fmf�8��(b�=�=��I�����\����s��F[P�# z���S6����p�B���������|����dN�x�v�݌eX��J̉�C3�ě79�GG��pm;��e"�����'��[�U8U6�o�;�t=#�}������ �Q�};g4T+N��c4O_��/�:ّD0����/�-��˯6��1<���d)#���[�ck�|����"FJ���
e�3�qͳf����+�VY�Ӆ%GH��g��`�
Q�9�X�ҹ��L&w�"�;�6�P�k�M���P"�{�߽ �0W�	zٝI�|Og?ݍ��h�1��F�>p�@O�5���V�;}:��0o&������){˞�"�.�{���bj�Xe��9/���1w?B�Ez@�NЉ
6^��:�w�!YR
�ߜTf�R�e�+sSVT|3���S�1ʺ�`�nzO_?`<��΃���m6��?�E�}�5�Oz}�{z�-uW���hImV�_]�샇ȝ��ll}O��E5�9�8�g(��G~~A����	�-�(�V)`p����g�JF��{�|�q��|�������� �YUP����yj�޹��4���^�=�u��{���ի�t�[*�^����� #��eru�p����ڞ��\�B?ZY&��e�〤ܧ�t��j�v���Z�$��_��Rq�WO��ߒ �*�����0��*E�K��!��WC{Q	��HO�-hlk]�5T�2���6���x��-��zl:KvkKü&}��c���D��s���C	��F�x��GU"C��P�M�t��8�Ҋ�N0oz���C:��7�?Aw��(qp �R*�8�
��=��{��:�r� ~���n��-�N�5��B	:N5Z�n�O�x���>����
��r�V/����б/�k_�G=N�`�"	��4,>��H��)���pg�K�ᲆ�����nx�@O~��>oί�_\#q�L>{|��kWA�����J>�䅘�V=���r�۵�+8���G��H����.�D;��cJ��i�&
S��>99���WA+��a�cn�ﾢe2��3�BX��&���Ҡ��L�ׯt8��w����� n��.��oh�=ǫӘ�F�$h0V-��+���������(�B��`qYgSh�}�<�����Bۭ%z"���bX=��������d�rL�%��);++fC��������PYM0�g���Ԛ+}����U=c7|IHH`��U-�wUȄGX�>=�8/qm���p��`�����&?U��[�oH?ϝ�h�Kx����uXP�ݛ��fu�f0���/%6��a&1 �C�ۆ��wmb����=��b�۳g�XAg_>h�dP�)W���e<�@�������܇G��S�s�����l���|��ys��f�%��mu [b�^�ŉ:~��i�?�ljk%bz�
j�,�֧�o	�:�֤�O���� 3a��Q��$\M�S$�D��[iXC��7><=����Y1ݭw�hi����Ʋ-ʷ*`�A��;�?xɶ�����8�3�7� K�B��+g�b�҅n6vK�!�<Py�Er��.Z�tg=�u��l�p��(cF479�ea�i��g�|B�<�����������I8<�B ����99�2��5��]�e��.�2��~���r^2BKӨ!��9��g�}|�8_����+]Q� ��9M��"�7���<Ck��t��FS3�j�ߔ������/$��30��x`����D
���<B�Z������V��Ʀ�{N�dC~�x���lgĄ���]P¯���u�E��Z�o�
�
�9��F{.�X��3V�1�׮d��v�eDr����1Ň�Pv�*����߽|T|u6E�_�gS�T�:��bz�(N������ɻ{S����7��-
�0f��y�l\-j��#wE�{�:�G+��;e��E �+Es>����_�䉗�ǿ(P�l	� �j�*�/=7`����o��z�R��S.:�r��Ux���_��`����%�����K	�)0W�w��W�g		GJ�}L��L�I��N� ��<��sf�� �[�R����qʅy�2e�劄F&��Om���eݮEQ���u�@����O���Q_�l�)
�g_����|MDv�to/�8�_�<�A��%8OM6���� i�k{y-��o���@��Z��n�?>;t�yFA4)���;㿛�5�~fa��ipgcj��:2�R?�B�(�Q ����������<=E��6=�B���)'�/ zSS_��e���oy�L6��A��3��Mn6���xD`Jny�'��Q�/g�d)��o���\��+����b�ws�y��H?`��AS.|n0#�NL<���bF��.��U��0��KY�Y�d����&�n���;2�!�r�����0[+4�*t�
+�W���\5�?� �c@+G	�e"�@z�XS}���1bڑ�7��<�-彺<t�9[S��$HyjQo�ɗ�.�x���K�.�>�@�0�����ou�0  �VlQplՙj=X-v.s12SW�Z��!9�!dj����o-@$�����A�=���ܞ���C����nM���p�m��Vg��/ˉ�_��Lp�����!R;Y#�ts�&� ,��m��JluT��AR�]�X�����3���/�	��ζ�P�3H��PeJ�uζ�ӧ�� k�,��	T�@zeL����%�B�Fg�[}"���)5���E���ȵd�� ��tY{�������MO�{(��)��H���C�f@�>���#�/�"�
�h?���"풠�5(,4;��b���Q���?�uI0�9LI�	����rGc��Z�$ ���%�E�S��bM��������=���>2���"45A�J�#J��Z6�\c+�Z�|��^��a6�7�9�Z��߀�zh�]��W�@�O�}����e`x��N�E�,���Hn`�:��.>�ɏm��UY�[7�.e��S&�U�a
l˘q�?b~�{���5�wiy�)��Z��'6���bbM;��^�?��m�{��C��o��K`{�t���$��q���'�o�y�E�Qgi�i���>�a�b7����5_EEf<>�Sлn�=��c�xmԠs�_��xn�Bg�����m��9��Tw����d�t�#����L���o3�(���SHTKds����s��o��n2�N(t4a���y�Rg���(�DAuOϦ��ԯ�l�J(]�@�zYII�T��O�f�"���^:���'H�� �����ҟ:O)W�%��0��J�+���/�"��ᩆ?y����U�(N�L���䤵��]�Ԁ��B�Ϋ�2�QU���N�n����
�CM1�nh�yʯ@LK*%:��w�J?+>8r8;]6��+̉���
],D�+~U�aץ��Tq'(}�2��sΗ��V�����E&�/%���HQ$0��3�2�0E����Z��߹�� Χ?>=���	G�� �^9����@A��T*���<�����[i��N}�ME��������ڋ�H�+����Yq9+�������Qg��7�rP/@B��WP� �K`"�D8��}��j2�'������cx�?G(s�%]��uF�m�߁��CPV�5(���F��4����y�w��Ґ���=�%i�^�Қ?��˨��aa�u��;#�����ө�6l��k_~b��o:���N��2��Kh�8;]!.��kW���<��&K����d��ol��Y������L��ZSb�'��F�2�h�����33)c�����|C��L
�o ]}V�q��M7l�����yk���o�yV�,M��Y�M�\X�4ppĭ;����]��� �m�!��*0����Q_G���a��E"��֕�}wm�����ė�f�X�oF����u�_g.��HLJ�P� 9n&��Omy��RJB�̳��Q����A���Sg{�C��#��A}Ǚ�>M��J(�e]��{�����;N��l�\c$�]��b��c�(��?դd��
��nݣ_?�1y{M)�F�^,��ʂ��K5~Ʀ�	�!���Q��$[+�E�e��x���*��n�	��T}iiJ-A����fg��o���/�N`>Gg�=���ӳ��g,Єfn�ZO~��o�}����? ���z�Зb�+N��Zx��`6ByIYR�?�p�� �h�P�4�/g�m�EJ%�.���<S03f�k�D�OG�q��򱎈���CS��/��xa�]���s"/�;<�<��6���fe�j��#1 �S�II�+�2�9A��z@�X��/yi��4j�p����NB�\��S�D��k��*� l[�߰���Ï`�e<ut�d��{g:<� ��UX;������'.[�I�K˿`���Vg'�ԖWQ�az�=�[\L���3��ou9�n�J��}`�_[vdH�7*���qw��k_�P����IM�{#��L���B�4ہ�˓NLe%^����W�-5������:vw�r�i�yA��.���{7�M�N���~�w�o�
p]������K��P_��|���6=�����s6?,����,ޚӰd����*-c���(rFZ���U���N�����ላP�)���0��!��rCX����1�(%G���g{D�����f�fF� ���F5rbH/Y}{��fcX��j(��x9�03�\��oL�?�g�ȭ��ѹ�ա�*���>����x�ԪE %�sfֲ��|c|�Է�&����HyӈN���>�ۖ㘺Øz��i�~�b"b[@p:3k�K+ ��JT�����wQ-2m�"���g�����9��g��F�G�����V<\�;�ʊ���H����Ր��'9-&\!���8�[�Ft�U0��D�}2�I�bc_�?�%w��7������%�W��!te�����Ý�`�}Tv��@�Kee"讞-�pn���F�q�Ag*��%���T��ѻ�%�z@�nq	%-����'r+�îO����8�X��Z44��7Xc`��ŉl��\��N�{ދ]�w2>1��wW �9����&&��Cx�!*����~�m.��=R `��=\�W*�j�}�c	��22����#&	���")�Fݵ7��� �0D+�������A(�)��"�������t���E���m�9�w,��$�:���#��M��i�y�4g�� �)�x���ra=� .\n���H�brr�]��:U���^.BMr�={��LD�'���֏��~��>���ںH�=�%^?C��U羺�J�J�4��X-o���&�-a�S^�qyG�r� o��U8(9ygz����t��A�<^�o+���~ �h� )�nV�����{z
WcҲI$@\>��&P�r�ZLlxF�w�30� Nr�E0@�Q��8/��3ߨ�_U�6�P}�ʊPO�'�c�$EEl[R�IG�Ԟ��\�G �	�M�0g~������tĒ��	3�4~�]��%T\�\[[BC�SQ�<� ]K��n�)/�
���5l�hT`m�?T�@ ��>�O����q���b'� ��Zv�#n�̌_F6E�H˪�~*x��߽a
�76|����� ���ٙ��+E��0��{==�w�J���B��6uc	o�;~��Y�蓰�ܜPK�nc=eO.8�n㮝��� �j�	�g��61q���S�Q�M޴q��Mx���*�W���. q���V���,��?����xy+�#Cԭ� R�3���ƹ�&'6c����a��Ҡz9َF��,-�����[��6������3u�Q~��Ri��:آL����a�3�D`�w���-���/�es�Os.F�YM�_��`�ژVJjjʮ�;�KX���U�X�y�EYVߨ��ӧ���`��~xϷ�"NGd��r��V;V��eώyf�,?�r�����jθgE�4��60h�ihX�˟Ů�<k��QSC%6P��ڴy����T{;�#�y���J�ӧm@�L�
�P%��h#GU���@C���^���(�+��x3��x F(�|g�D�&�;4�����Ol@�ژY, ���?����3{D�����+�!!F���Cz�m�L�8R�X3�ﱈ�_�'r�K�6N�q)<�efU༢�K��Oҙ P^�˜k����N��g� q�-��7of��Q^��{1���3����huqqs{r'R��T����5Wx��Bs�[8 J	��M������ǁ��Ύ�%���gϘ�n�L���VP~���W�+���U]�;�}=fqW��Q��Z��&���(-���-��"�#d�:[Բ�PR�J��l-?�VOF����t[�"��V�qY݀��D"'s��T۳A�>q}SS8� Gd�o���a�zS��c�D��NSS�Q-QSK��M54H����h(�e����햔:�QK��[�Y���.��Iʞ�rS��HK(-.ݨ���5� +��1eG%&����IK�{:��\]�+�?{uIw)X0��$�|Vt5/osK���+M��sdFq���sע� ��e9����d5��F霼��Rū#T��U����hb�ײӦ�aiU\\���s��C���q?ƿ8���1���-����)滛"=YY��2j��y��"��j�%ݜ.�3�'�4r��� ۝<DG++��gL��\]Ӑ�{��?�x�7�A� Ô��Êv�t�;;\H]��[�^_�������\�w7�ݽ;����I�y�($�8�ˠ��ǎ���Ϙ�q>�+���&�l�:u*W�ԁɅ)�XZ�Gӊ���hb�Y��zcs0�P���G";���8;�Vդ�[��Xpw���:���"]W�9����:a��yOC[Gf 0I�p��3�ᳳ."2ȧ�:Q@���x �'����H��+��&��1W���3L�'`�J�]*jmhx��7K\m���8��ZZ&����XYv�!�g��:�,]D�������C	�\��V��('�:zD��bz�l��j\VցD�DyR-6�jxT��zd�`��,�lm}��^dhh$�k?C�Smh����S���w����/7T�YE�r{*�? �a��:������i�.��z�N�LaF�P�Hg��?XGq����mxex:��%���33��x,�{u�<�R2]qeM�r��z����Q��E�`����"Q�V��4�/_�~��?���
����g�05��o=��ػ|p~ߺj�<�`L�����a_��z��Ƶ�f,��E<�%׿&����>�_$44(ܢ��1�T)��$�Dk4�X�.x$��Еb'|98��4�L'+��ϟ�%&�����$#������#� ϒC�ߟ�Խ(�0�s�r�h��W}�I�3�R{Ȯ��j���OK<b��	�'Z1�.�n�E3������!������|aAƊZ\xCOIT�p}UC?R������o��H����(T��#�m��}�T���i�W��1Pkt�"XMc��~���ʽE_{�*du��T؇��Fk7T׊1�ǖ�L�0}�ç�~��3��b�%{��!�,��yr�$�1����Su�u�U%��v����Y�o���}������*@�!<�jP��R�=���!�;!y���`F�o��նr�f�~=]��>�Y�c%�Q�bK��K�>���.��RD�t9�k�\��{�M4ΞF��<�H~�P鏉��h��k��Ϝ�z^���U���q:*Z\yچ�z�gzh{�C�[����޺�램��� ���i��y��**�����P�Oc�!��q)�{P}��>~��q�ܢ�U	�|��C����Đ&jB����w����.M�0�I|�9��b�[� [�gOk�/N8��p�v���`"�$D���҈�X�П[�Rƌ�ש #�?mja��]�j����@%]���߭�yP�g�3|�]+c�MA�A�ꡖ����iS����`��\�ę=�w�y��؏�*�T�u�Z�����U�ɑ���k��W�=����J��[���󈐀-���m�(�2�Z�x,�r���渹K
3����7�O�s�b�'-E�Yn(��|��_�ǵ�Ja��n��ǵH�i0��kt�JM�����
s����'��8�?[���k��v^��v������;������;������;�_������5	|�a�
���;��؏�[?�~l���E��ߏ���'�~l�����c��֏�[?�~l�����c��֏��/�.{,�����+�n���h�N\=�W�	׋1�1�
��xo&P�\���<TQ&Y�q"Ź/��ގMH��R�;iy��������˿~������N��O�Z�����1fj�]�4�-�+�k���L�a��I��]���n�B��������^�+���m���BߏS��������){]З�U�|�Y����7zz��꼨��Y��=�)�Yk��?}M�jk�a��S)B����s���������tA��*
}%���t�@õ�9�񋰽�,4):3B�*J`���B��e6�A��o6�o����k�.	��D���q}�������>���o��M����.n��+��8r�[�����.�yM���|�C�?<��}�qrq ��7��/�m
}�:n���̌��o�µ���T� C���IP�١\*4�ۥ��4�b���Ŧ�h�>��p�FA�����;ڧ�//]����tH.n����Q�O���E��[4:>�/�}ʇ�����@8��M�Pl��� �4�$������U�]�y�A߬p�ɑ����B�{JEK.�߾������LE	�7%lV7'����τKF�u�߰�y�;�d���z�ף㟣�V*q��/)��I��Z$��צ����C�B�����C���!�_@5���(W��(���v�Y���\��k��Y�i%�hx�r�?���e-V��S�8lv�\^t�W֣���|�.Q���#���@Ay�?v�e���VrBo�	�������YJ����Q~ڠz+Ep���;u%����;ڿI?��B�9q�M�+��4�O�(��ۂ�d�v71�g`�9H\Rcww��t����971��ndd$�C�o��7(+)q��⳱o�I��#��!VI��v%� ��1@����=�"**� d��e��"�ww=�+�]O��@�K�8��^�.P��f9tO�f�7�:W_,j�����C*����q����PY�}ee�%���;��u��e��OPS��0�L��6t�2�!�Ԋ�	�J�eqǑj�`��������M��	fbb�8)@P�p'��\�kI�G�D�8M]��4W�7�u-���� _[��g&*�nD�Z �С�Y��X��ᒀ��9o~$@K��S�FPj�7Pm��_�H��C��\X5�+�{�5�!ǵ1ƸlA`�����̲\TM��h�m�"�g ��`%��*����b��am)Z��ԑU��h;8�-类;��B��uG�T�J�`��1�a���v(��t|���V�'wwu%�(2QQ�	8x��M�]!��G��X�!��̃�ammmVV���Co~���  ��'Z���kӔp�ySllk?ӆ�?U�#᜸�?�`�M�---=�d���eg�/FO��srh�A'�?:�0=M�*��P�]�"� �ꈟ%09���T�R��M$w�|��&����C�$p��E�V�"�˰�K�vF�Z}O(V��ZN�е_ @z��J��<���~<�팘�~wR0d|G��ˍ�I���\�X�w��f`�SR�H�4�ae6iu� `���LNFX�p)B�q��8me�������ɷ}�`àOܭ�Oc����u�;ݎ^P�+{�1r�4����x��R�e=Dˮ��~@� R�;�ӑ�Km���ߎ�y�ǓQs�+�oBrr:2c���gԔ�$=�����-�.� *��/��P��Cm�8�����B���?c3����I��$��B���� T�6k
��Xv�@�P�^M�:m-.*�HPv��}�\Hs�A�ǀR��yH�� ;� ��"PR�R;:/�z�j�#��`o��	L�MR��?��p���S,����.F�r�p "�r�ɣc�b��b��N�-�'��GZ�w�h\T:�Z-�vy���G�V@E����)�wtv2�.1�j=�zn�)�/]����W�ĸ���v/{��2�̓71�����UU���j���l&EEyD�$�=B��� Q���#ge�+P2�1���=�	���Afi�8( �p��0P��%�Rڱt�g&���Ƶ�}TO���B郻��I�'��E8 ����mc8P�:7A��^��n~��ys�m�)Z�|R�yX��sH���K �� �')U:�<L��y��0��yj �C�2����b  K�{3)rEE��9!^8�r���k
gAX���J���f{ĕ_�컀�C}F����&��*�*�Y-�l�*�hY~mHNN>��Zh���#��azT��V`*ճS�h �E��������Ǭ�0Y��� y��׸pv@���U��tP��g:�JKcc#[F����815W]�CՏ��*F��h)����g�T�$��
���Gb�:v0�p`̗��!`�\>�.@����L���[���� <fa�<OL��֦X�q�[@�ٌ��1�Ud������Gd�����Ǘ�&
8n[����EnJ��{v�6���	ǌ2T���A��3ZUV��0>��z���<� .aąs��93:
A��:�D�޻�	�7T,��Mb�\\!vh�|��)��������J�j���R�`�TY�(Dl��\��@Ԋ"�첷V��P5
B ���,.,���1(����Md�fNr/���?��9sf��yfι7�l�w������..uW�Ӛ�Q/Q�����u
�4���yw����:��r&�OS�B�:K ZG�3	LC�c��(A%#�M�T�pG�a߻�fӰ�e{$�~[J$��эw34��'��\2�/�d�OԾޢ;]UXs�x7�j'��-�8a�!�w�}�V�ߕ���?e<;D^a�\汳��> ��j��3��O��`)��}�١�|9
j`��N��)���7��9@�f���`^yY����WhlM�&P��'C�jzw�H}9����w���9(�Jm�#>��&�߹��G�-	�-n�6֖���4=Id8��f�~��c� �u�x�<sΉ<mA�:K��[?ɉV������i�R,��5&���$�DSe�YIKe��1��`��u0�qǿÔ��2�!�q~u1����n�A�xa]�%�Yi���D(3uJ(���_��16�i^,�6��v!8�'�el��$?�)�QHXN"U���DW�#��Í(S0��[wz�����ˣE��d�4��Ӣ
=���O�}R��*�}q��I�o��(T���zZ��)�7���95������w�/ 
||�c�k�J�3���b3���p������R�c�w˥�͡��wi��T�cPo�|���`�zT��vH����x�wO.��n��2�ǒ������\qy���3�W!�m� �Rh����@�]~2eTT����0_*5���nB��[˲;��(p���~� ��c�_W �E*��E��2e�W���ڰ�
)��z�ѥ��̢i����
K&�<���v���nkg�%���\�%~i���B�&&��A�y�D��TŹ��սc�"CD��[�0
B�)O��o*�}U�ݺ������2)4*J��x,&L�qGam��/8�Z�6D�oPk�=��!���<y�$(f� f*z+D�����HR.g\����m� ��<�,0hEzMލ�ք�d��x�rf��4.Z�F~�K�+��H׼�81��]a�oE�v��G6����'L����e�T��>���N&�i�5����6*���h�y��w��#�^����.q6E�Zq�_ډY�݊�y����5�&[�����`-���_Q���k���E��]�Zρj��]��={��5$�S6�d9�o8�ϝ�s��z�m�?��pn%�ХH3뚛�k�<=,��>��R�c�����
=?��DD�{�מ���2p����)��@=^�y-��>ҁ��{��3(�����
[�M��y/�K��j�;P@�"������Ԯ�\�Ө^ZX5�t��"7���V�e�ye�l���?*T`�l�D�3���.R�� '�.T�3������_PK�C�{�Z5�{�H��gKK�W�P=�/�۸�8^������%zz��I�Ĩ��]�($_���8�Z�L�$��c���J����T�[ePA�W�-n����i���m�YMt��I_�@�h荨b��҇p~�ܨS��䘥�U6l����DS��!//��I��d�T�*�z�Qcwp�p'm,���-�I	�5�F�k;���v�Ռ�u�?�ZRS6t@��+��%}K̻��3�+"㙪�S���Kz� uv����A�l2�q�בV��<��dk��z9L�Z�
'�n�R���b�4�w� 1)��rp����gz=�?IzO�f�]o޼9XS]=C�`��=���C�1��B1M���׹��5\���'_w�b]o���I~5j�t׫��P��u�\ۼM��(USv�p��p��P:���{E�w�׉�r,�78<�y���i
����Q�\��&��+��`�IB�u�hx+���_�����eb9���'�QķG��wqr?cD��Hz>%:5�`�0���ҝ{�t}U�D~��7����	�gɦf*ԸK��Hw� ������_�>gK���^3a�u3v�,p�h'�x��J�H��aN���s���������lIp����)֥�pmF�E�����$4_Y�Xߒ���Ιk�Ԗ^?�e��`5[m�$��)ƊL�"�Ҁ�����89�e�y���X`kY
_>s�����'�Η�c��}6�}b� iU"�Rm¥�Ӈ7�Z��N��}�.ni�E.����[�,;�ߍ��]��<�c9�!�Y)��8�Y����$�h������H��K�4}iU�Y��@�tॏ��Y�9/�8l�x�m2�]���Q'0��V��?�1μ�>�A�;�dȰ,��H�i�ĸ�E��^l��
d����o=^��-�x��	n�O"�������M�F�6v籃�mR����(����!�W�T-f�3㵼��bK����))����E��%دcc	Z<uh5��"��\��s�=	<.��J�������C��į�Q�L���c�!���B��jL�w�<L������X�$��5+It*�����'��LU��� �P�4�P��T�"��������q��I��h�8ހ��c�C?Ț8P�
�$b�2���<�V��S:8z�'�u�H�l�_X�o_�4���?Y���{��s��7�gXֿ�b���{YE���߮NO[Z}��__��u��k�������W�t��/�}~�r=�.�L�c�qo+?�*è�Vm�ќ"���Qmc���_+@V���]O�
7��}���i��ɓ'�$�i�:EfO�BG�y5'�[���wg�tΘ8~�b�=.ەi�~X�g
�K�a<��d���p����P��WۮA��3���jhd[�#t��-;������{�"��[_<��\~��օ*eKa>�$�$"�G�)NH(8<?M�H>����4�./��H=���7���t�yc�#!hU�i�����[�N4?�w��؅n'zӷ��v�-;Ў�AP�w=7�KGy�)�����x����H.WhAƪ�(~����F	b�ɅB��O�#J^Ң�$���P��A�nQ�-�����"��ϧ۴���~���7�\S�Qk���ؒ��F[H�O�[�`w��fO��zG{ޥa�)�l|��Q�l5�竅D4�"
�{��ʤ��?p��W�,Y�`�<��1����\nQc�!ˍ�z57��-Mt�_O|w��rc�Н����"�kɳ8��������(T�⤶ƢQ?O�٤1[�}1��9b������L�|����������}~V���Jr��+[����-Q�J�vg%:i�#1cTQw1F����0��� gWȒ�---}iJB�_�mHN6fv>���gXT�co�=٩BgM�=�Bg������Z��l�AvM�y�ۤVG��p�� 2��w�L)'�b!q��J9�� /�]�h �y��
�z˥�ÞQg�ImO�Ԭ*QC��}:O�(A�+0��������M�J�f.�!L����O�0�ߝ�ȑ����*<����AuuujP�9X�^ÞQ�Gb=���h4����>cSJoa�S�2���B�z˪"�������lkW���6(�V��0�w�z�č|�ԙ�o�O':��)b6���8�F���-8L$��6ZV��SF��@Ss؇;d�>|�pgHȈ^�*��3��*���ǎ��Jf�������J���s">��(l�Bh��_�t���C��)$x�Q/�^7٤��m{�YfW����:v�<��==B؈���|�Z��|�L��,-3�B�p]DP.*�kw;���s �MzxyQ7�Т�Q(�F^�d�����k&�=�e���\[�����k���]ޕP��N��W�������G�[����j��A���+E��|���~X�@��8���L7�����ۥ0b�
��w����"Cm�w7T�I|~I��gݻ�Oij�Dyo�E��?�5�)�h>��kd2�������i�iɻ�H�xy�����s��
GmqQ�o@ na��� �L���_��u\xO��ΓJ,���y�u_����5f:��5nٝ�b��'!B�Pa4Al[CA [�s�l��GfĮR>j��(�0S�]͊E��ڥ >1-
�יe
�?5�w�fGp�ߨgv�It�%�,Up�����B#-�<t��s��?>o�w2g�H��82�/��v�^�E�Hff��$uá�D!O�R
٨�#���dN�	�yCh���a�}����F��J�1�F���y��Z�p��I�����W��[���۲��݇��B2�<#P�w���O���ų^!�v5F	��)�1���ʸĜ��ڀ��;�Mir�Z<1����������s��c����ξ��J���<(z�B��)M�1d�k��u��������I�tY��޼��?��#�>&�`^��"�����+dwhF��{�5(�-���P��{ o�II�ƶb� n�N�-�R7�����N�vVjʶ3P��L�(�Rw7B�@��G,�R��J��T�vR^ug���ѣ� ٜ��Go�Ȣ�޻w�Y�;��MwJ��4�b���No-O�wk�S�G�9����9�L�:/
s!���w�.�~Se�hNg~�)>�ȂL|�Ν;��z�6
�)��%��f5OA�S'7>��QFB�E���4.��aN�?q��?7��tM=� ����V/�	z��"~n~Zk
E0���@��R��F�w(Jk�����J�MP������)%S���i_�Oi#�`��	�2<��n��^���0ϙK_î/��zK�WG�2)
��C�ū#oƐ2G���3�����������\!�+A��S�%'��L).�ް�s[��nS:2<8:[�3�Lff �0�ܲ�����F�w83�u ܘ�%����Bn��u���Nl�
6Q*�I�n�r�װ��ԝ^�P��bD�R��?��s����� �`��@8|�[���(�LE֯3CGG��sFW��8��fܺ�Z1��}�@]� bX���G�{	s����2����K�9�(��F���{z��$x9�A�6�T��+n^�}���g4��9�k���Z	6�:���DR����{�i�&�,�Ǯ������|f�)�������J��k���v������hcJ/� ����:@ �qM6��" (Fg�X�{x=�ŏX�v9��
�b?S��� �L���H6�a2A@�,�&�b#��
)kZ���!r:�9���l^���j����H�#�Ϗ��n*�P�u�'��J&gj�������^	[C]��X ��|��<U&����D\s6���~M�dB���#�}ɑ%eն���4�6%Z��0џ)MR�?/��[E�*��O@/�k|�%��s)LW&)�Zka�ZY��j(�] �;qK�?G�l�k�!cѫ_���5���<�q5�)s���d�\��=��-�1��]MԼ��Q��\}�5x����P�&�υ�VO|�_N.��_'1�'?���X��iS~Dx�tt�b>� ����Eɕ-C��1JO}ww���aP�5Bé.]��z��l;;b��n`샱�7�֧��G=#�����A�Uٙ�oĝ��G�'&֢L|����Os��*�W��v[�:S[?���N݁����v54\�)T��ׄ)�������BC�@�����b�0����=SA��h/D��Ľ��Ə+�M�i���9����[&v��}x�#ۈ�ϙ/4�(hx!� GK�^�,��m��0�.��OtvvN�b�/�8%����]��,Gi������@_^�v"��555�j�N&%K�%_�O�$j����qI�R۞��Vc��d.��R�;(��i&%	�o���q��IwB43�Y-��MgFa	�g����N�9�	���$�a��
�F6sU�=�SZ�Ty�=���<�p�I~i�o{�n~"��P"JKk�t�`�EI�C����Z?��� _���?F����@F|��-��"�\'��%m����9��ߺu+��0��oi
�6B��_M�I $������3�~
A|rg�7mU�1~�����0\��$	�n�on��s���7 �����f�
ןFk�0��RB�pB-�٘āOıwRO	��P��%�%Vp���ɆҨ��ɅR��Br�^K�Fs���-�w׎�wS�;��-���4�73��)n�LOq�KS|�mo��#��"��%$aL�1>/J��k�����z䓡[G'����y���3�/����h���_-n�ĴM�9�52"�+�/���e�i�0G}[Pw���5iiD5v�(����p�h;G�4�o��rVH^Ւ�$X𲡸4!9��S�����i?�J>�`%�x�L\�:u���qS-Ε���m����>l�����Z�Qw2�����Y�a�"}��2Hm)��n_��If�C>m|-N @�! ��Yi�1o�[3)'���6�Ό���H�풉C��bn��(�S�l�6��ajL?�dS���s)9�m|�Mu�|��w�K;pQ,'I�=�ԩ!c܀���x���+[b�힦E k�@��Χ*�"�N�����3�� ls�dq~�o�U"�v<���z����e��L[u)��
�4骵�:�;sq�VNS���ýGz�e`��uF+;R��?inn����÷�l��M���JNA�i��Q����?��>5�y	?0Ց9,5���լc��fz���WEE�qS]����:�+��Bф��&YB��q��PU{�{�^o&k/���.�l	�͊��y���\�5#�$#h���a�?B���'��&�����Cjb���s
��7�=䌨�A"
 B�E[�Rq���l�N(�Ĕ�B�dh���S/<�Gaů��v�&�&p�t��"��N����fH/��	�R��g��<c��1��0DކA�̉��c�|�8����Y;8�ػw�I�w��Wf���5P!b�f�۽�L�V���B>o�O �lV��.�{kJUn�SL��>�C(8�@K�M����K枕h��-C���XE褛?�9k--[������b'��L YO����|K�р�C;%��$���$`�v5嚸z8u�A�Mm��{���=�nu�'�D�&%>`���J�����ԏ�;*��|Α�,6�$H��S4��{4iۤV[���	pxlY����|�xj�K���+��3ձ�W|�x����d+��r�gX��ˆ��a���/l�F���|�B���#�P�Bv}�p�����-O���[Ba�*;��0`��=���7�ŷRU�z�z��I��s
�W~:6yv��[0kͣr[��6�-9"o�0�z���:��G#���T[B�*��#�SZ>Y����s���K�b&�춃�Ozc�C?��N�h�pܫ��0rēA��a���6~ˌ�r�Ġ�;��GIc�4��Rq$��#B	z�K�J�^����
�d^�d��ifl��d�L=��tBXۨ����ͭҁ��Q	q� �J�u�]�B�kN����,rP��[�����I�O�h���M��`��/ ^>���֒0=H�bQ*p�]�-x�f�,�+�®F����dj�D��3�v������π�+��Y�=�{�����D�3=�5��B&�\Q�	�>��$ޮd�O�J2�b��iK�o�,�N��e�}�W�)7W���g����)��׵���kB�4f�x���.���$'_��Ѳ�^�{um�y}�:�J���F�P=hM/*�CS�S�|}��1,��+��m�"Ɂl�×�@�mL1@[&xI�I:O��n{zE�Y}C]�9��j�������li�7/؈�?a��[��=X��G�)t�*����#$J>�"��/هz�C�����.y���7�=]�3�ض�\i�W߫B:Ŷ� 5��8�oyb�l�7T6YY�[#��_Lɲ�wa���1#��~�z4��#k�/�B�%�Λ������P@�`:��sێ���9�U�h-��
�f*��s���PX�Z?��P����ɌMh��$�K.�����'��bz�zrO0/ �]�vͮ�g8H���b-�#h�˩�P<�dسK7w/���J���U��!���+kb?���\�$"h�h
)�.{��9_�^8��K����9w�x}�����O���̓�-�P�7��}Y6��V�6��7�~��w�p��`�Q�<9��IĤ��$�PW~��ݯ
�g�G�>���H�ܑ�hg
~�+�k��2�&���[�6��_a�ap��S[':n|>�M�-oFۙ��"Uf	j�WB�8�cJ�L����kZ3��1��A2�2�s�W� �� 6�z�fiE�͉��e��,�#_a����Ȏh4�N����ѣ��e�T���%�=�0�ҕzK�4,V��N���)�b+��D�W>^�ũ	ƪ����xH��	
n,���xw&Q��l�B�F#��^���-P�O��oM��.�+�ܕi�.R�I؃�t�;�%�$Bu�����YR�^�2�О���@wz���!��<{�<v��t������.n
��G
��^r��cK�ÅE0-�	����Q��Q���i_vm�\��0z<�����9��&`�{Xe/SSSup�u��XA�%�ʕ.{4��e�)���eo�ī2���{�ؾ�e=D���)�	M�zܡl�[U�.ǀ	^=�T�|� �eS
�s�@��	�1�N��ìq�:��-Abc�z#�jv�������y~E;!�_Dl�S'a__��WS]=U���\������hkkc�Ǒ����d�Fë�]�H�+��>|X�Qei�0�����M�Q #S,�m�YV�n�,��Fq�[�O�5ڃ-�k��zȩ���y���^��:Z[@��wߔ/_�ͫ��O�շQ�c�ՓwI�yC�ȼB>#�w�<�传�w��)j�ͻ-����\���u��B���������P��W���R��F���?��7Ae�h�����%}p�ZM�Pi�Sւa���k8, ��z��*K���Hl�-1F����Ta������*���-`�y�M�x���vÅ����n�\y�'�ƿ�fa?^�~����]=��d*���rb�k&8�W2܁>gsK�L�y(&ѩ0��6����x�O^���d�t@�s<���1�5BuY��E�q)�k��=d�z�F(0�:
�I���@'?逦��9qѣW����y��m�+�H��)�,f�6	fv�S�Q��ᐢ�G���;�r���[4(^����I��9N�3|���f�1���+�1^l��[�W_U����vZ��-.NW�{%Wzi-k��+����J�&W�������w�)}{c���7_ٝ]�W��{��O|��-��EM����}�hZ[�Z�� ��s����t�\.׮�[2ͤ��s�{kϑ�iji��`�\B��#��o^Q�W�/W��)��y�!�(��H�F�Pb��MK7g/�	�/�a�pϓ'Oҁ�����ȣ!r��h����;{P}���ȘD��s����p���	}�;SzX�M6)n���É�NY$0�Rm�b�w�K��U.�.�����e���?c�|P͔�Xwi``������e�
bŃ��-�Z����@)�Ng�2���:����x"f���h�$�Ň(�k���ů�n�['�����Ǐ��kɄ�+T3�&A�>'�"}�`�̾�q�
3��2J9�s�]���cW4O�O�n��_��;��e"�gZw%i���Dۈ����I�j��"�Gݻܐ�esYD�K��| R�%�vQ�����Oâ���l��}7��?��G��O�v"� ���2�HF���ħnj��r�Dۇ�Qq�8�b����O3���;���԰%���,����LOK3��e���a����m�ήtw�qLF��2����C^O2)9H��y:>�p�L��dq;Հ��,�K��ˏ
�m�%!�+CE���)�\l���7�K�d���%IhMJ��2��$nn��+/�t�nS�D�	��}��>*�VBIfWc�m��B�y�l�}��~�ŒU��V�/V3�S�-���� F,'��+z�KK&F�B�m�<R�dxܺ'��(��"lD�o�*�qb|���
���hk��0�]��Y��`K��ml�#��Oe�L ��Ni� 2��/���ܼ��ſS�L���Ȇ��
���6�5�N�!kS������r[�*Q'�t���Z{?�5��R�{Xx�I~n>��gI�U���s�2t+�q�J�}n��Lt%F�P迣�1t����-+%����<�y��$x��0i���GK��a�l�_���WX�S�Mg[�`���i�]nJ�Y+ Ch%gѻ�D���C�&n��m��^.7������G�Oa`�[H�χ��vNR7��So�g�����*�l�ӣu��q/�̸� #�Y��{� �ߡ�7��ٴ��,�Ƒ�
gt�o@w�
&,Iu1�w���l��nZ�2_��A�"�!�|�:|>�FZ�IO��Z�~�?N��`�D�5֎�9�k1[��(*�>��/u��z�@+����Q���n}�h���Vd/ɢ�un�S�+����]E�q��k��a�k����bE-c�>L�:���t5;�:���^�w��<O�+�% ��Vd�c��7#}Q���R�Q5���o�BI�s�͔�!�v��ck"�1�-�v�q̬lɟ)���U��)�8�t���Üv�.��	~���s�4�[(����Ȳ;��t`DV֤�NMN1`�Og� gvF)=5UmW��)�՘��v����}w�Kj�
�x�tt<�r���Vt��	�Tb�&)su�<���D{���K�F0�"/)9�|^�	��2�f"��b��K�y�F��~|�~Qs��3tJw�z2�1E"Ga�V�/:J��PJd!�'��#E,��hG��!�~�Q�;������ %=8��\�%����*��VI�WVV��e�b*&	���շzJ�qK���Gijj.?�@�M��UM�mj�T\�d�[6�@���u3��"B�ڤ��)))I�J���%�Pe����=��:�g:�%x��w�����
�������ȓ(#���p���%
/5V����B�ק�R<y�^:
x�^�^���I�m�=[F]���֚{�3�	h��Sj
�.�*����)�0�XZB�;:��W��;���FԞj��6Z�6�|�}A�É��e��>�a�ǁ�����c�y�6�r{�n�ڥ-�)MR�E�C7��bF렶�𒪓�No�7^P��_�9#�!�~������Os}Z�k��v�� ����_�񸮮�!đ(/�o��Rw���WD�\G �����(�{�����[f�~/��^i�Mu-MMW���朲޲j��c�)�i� ���N>/����m��U��f�1�'�$j�K�4q�*c��`��-{�9I�I��ʀ R��O�}*�����KU�լ�lY���D�~OX�㟢�x�,--���s���~�U�kA��L�7C
��c{m�i~�w��Cn!)r	�8��gϞe��>����b9��r�,�Zc�Q�̶�/�Z�������﬑XV	3Y;��ބ\`�)�iRRC,x��S�w�1If�P Ly�3| ����@n/������xe���)�>���ݭ�]Ky��ƺ�ӧ�Y vz�W���
	9A�P#�A�Ѓ9@��{h���-tڱ��}�,����&n�ٚ�zrp1�����z_Z�U%R����I�ۏI<����]���LN�eItU�1;����ӧ7/@���%�I�}Nh&����hIͰ�*���?�5O\`h;�	�6����>��C���_p����H����*=���Oڢ�=\h5�x��	�?�*Lw�J���A����"�ҳ��һ��W�T�tu��s��/�<�����7�dK��d^����x��{�t�$�^J)Z��"2eK���Iyâv���T��G�����w�"��
ɥp�r DiG%[x���	��O�~*�％��qhѐ�~�wL#I&6�I��D��H�֯�Z��^����+>��wEid��̖���u��o�V_I�Ç�u-��'��.x�J\�?$3m$'�c#��W ����=�'3����99����t���PM�s�|�l$��͆-il�0�r/̖�ʲ*��yVs7"��^��4����YjH���8 ��!KEa�P�g>/��oP/�QeQ��+�}*���k#兑�,�����[�v3�m��r�����z��t���ׯ-�΢_�=�)�*9�>ګA�y��U����2���R�S�̄R�6�Bq��/q�94�ï�,�����2�ZEC�1,�ܧ�*�RgSJ�EaN!�W9�=i_�H@��tG�ֻ%Le����J�`o?��h9QJ�`N	�i^ҝ�J�s'�x��63���>v�סd����GF���'KD!EN1��:A�9e�e,-X�vr'��`�yqwh���N��tzN��v��1G�+Q'6H�Z��\ûh�ik}]�������*�Ϋ�o�B�v�B��sꀗ%L��I�\h�*���ak��Xc� J-̮�dM@�*�}��N�^e|�d�Z-,,d�_�Η,�0��:Ρ�	u����T�U�,�ws\���Ȩ���5>�D�Ә&D%ǒ(Y���dVٵs���wĹ���)
-"ϓ��Y	&�jw��@�>��Py��%$��]�~ɕ-A��݌�ɆHo�����.ج�!�zD�����Ѕ����{}p�y��ڝX��N7�����5����<�/٩G�M��dD�K�������/�|a=x�z>,A��l����g2י���ٳb��-��lTH���SKK�#�J�frV��\[H�D��MU�!i��nj��>[>�LM��Ԇ*�Ϲ*[��|�ߊ����{�����0_J��/����T[ufƆy�� \���3L`G�a�o��)Yr�oPt�`��=�r,0��ݳX��%g0.8>�}(�����n���z9/99M(L2)!��rU}yP��+�.i3f%'xI�T@�ܷ�0xP:K9L��9���ٵ�2�S��䔴rGw���*�cդiH.�>���~�.* ��H�FtI�����p�KLyN2p>'t�C�tl��j����z���NU��ʽk���G:�y�ƭd�B��K�C�� +}e�Q~FqbL\�]J��Y=�)���uq��9���4���eW=QDV2��jM۬-���cc���I�3�5	C���Y��S����ROi�Ye���ߌD�1���H��}"u�8���<�L�*)'3��(������ u��������ڎ�`�r��kkk��� �J�~�Q�qdA�x-�ɰ��:��n!MT܁c���������wB}�k�)Bs"�͂���^����ID�$Ok\�l^R�&;@���Ν5`�	�RR/����ͫ�F@Ѥ)��Iy�~e��*��%���3lQ�ѴvW�''�g57c{��)�7���83q-�l0�Q��F3�ڇ����Oi��p婴����swϴ���d�>/��Z��ݘ��ԡ#�1/�r`W��:2�:��ws�-�����Ɇ��X����[�D�Z��*�0����y�Gp�+�4��$=�)���~�����$B�3�eH�B������0Ԝ�M��B��k2�$�g�^fW!�Q�	>S��m���W�W� ��$>������>hb(O0�T%��%��=�3�����Ɛ�hC]Yh`�������4�)��|���m��Ii����E���yk��U���Y��H���=<ğ������yb��B�B�y�-�B�ZF��O~V��Q������*!'�w�} Q��	ޑ�1w��jFX3ԙ�İ�eG>��χ����C>ݝ	�E7�zDT�u��3[�H�b>R�
��1w�¶?Z�n���#��C��v���N^#���X�pA����:{�厴��6.IB��$:����<�L�Z6�'��i\B�K�JB]�,�jL�8|N56�@A���Ax����=��s݇��cS���k;��6YY��Z ��������0-Z�og��Cq7��k�Uq(�W�nT2f���۽���̮,����6�m؝�F�r�=�T���aNJlݟ�`H5��*�s�y��h(�F�Q���PP@����C?��MOi�۾����u���f�c[Yf.�5�A������G��<�~��߹��(��Ogs�sds555��Si4����M��i"��6)M��(����? a��0�lo����vt����|`6-�R����*TT��,h��C�v@��1�Iku&w�|�ip((�&��)t0��$�k�%���la�k�Î��K�2�W{�)&R=|e.xρc�e#�===��(k��u��o^(������tP����g||�?�kqT�}ܒ��m��Vp�����TQ�T_''�+g5�[�3Y�{����E�_�*cRr�&����%�r�ȧւ�I�p:���\��x?��Ǘ���u��yG��)~�牀y��<z,7��]W�����5"}|W���ں�-��*��[8�����5�3¿�;A1j<�ѱ��E����i>��k�tP�!�ʀ�.���Ӷ����������	M�
1ëX_��ЗDlkC�V�rZkQ����D���'���ebL_����7_oY5��܆���4��4<���� �Y��s:���]�K������k��o�U�Yv4B��ni��յ�1ޯs9�)%31<6b��&�.A�}�%i4����W�2M�NF��P��台�X�l�jV%<`�Ѡ?���<��s�Zn���������~�� ]�{1��hZjj�Ld:�٢��-!�����������|��BE2����3Sa:�!�z�z8�³5�E,��+l:���#H=:�IkzVe�福��x
���$Q�r|55�;��
�Hm�x�q���K��k̝�?GL�f��>w)?��95c٢E�9-�^6/BM}���e��w�Io��~~>��\M���KC\�٧n��8�=����e#������"��y�17 ?�_�~���5{y0p�'�4��q4$P�8�T�ꄃ�z�S�>���_C�p�t���t�UL�M<�3�Y�����.7�sFX_��liiI:1vj�P�`i�wb�1��<��kZ��C�w�eU��R|�Ӈnc�<A7�%>y�)��n�XOybH�����;+�j ��!��VA�jYN�����'>�\�s����Pt�c�6Ӣ�Xȷ��w{�\(�/�c\;(c������ҒٕZ,��;�[�0��G�%��D����OvgگǗw��*�~�)��p�_��[�C��*@&4��ݧ�A'�sbbb����k�ل�ߣ�`��i�.BhD|��h���#,�Ǝp�ִxO277_>�e��EY�#kO�������M��u�bSB&6�'#���R���TIg,[�Ty��ah|g?�2��HGG|�_�	���R|������ii�Ȳu8��昁ǂ��d5�8a/��!��8vj\�f�(l\mB/\��D�pb h��}�FwH�0��i���I������,�i�6!'�=_6dj^9��>D��YNn��<IO�P�@�d�ڬv쀎P3f��w�(p��jw��V���� �GֶۓN�8��Z��
�N�;��sxJ��'k%���C!k
�iI<�ÿ8��
8�n�R��ͫ��w���&%����%�˿7A�Pv�14�����/�{����IY�m[��U:�z�����7���w1Wk�¬�*,v�W�ε́g�.T8F}}�3%�~�u�p�x�������C���Z�̼��;�����㠾�Gy�95����/;��[��������~�e�n]@��4�j�������/�yٵ����y��w�ZeK�6��UP�?t�/޾;�MD"m�0'Z�~�e����T}����.�Y�Ź`kF)Xm��m��i]��+&q@��9�e'h+������u���RO�0��u��.W,`�^4z7fgg�U��U�h�=���7>�	�`%>�d�ȝ��3Fq3�M��Í��N��6�1�*������hS��-�;=.B��;�ᒖ���{��~�Ȱ���3��Uf�q�ƫ�� ���`�4%	���]����3)QB9U3�����E��U�����/��̄2�	K�k^�����J�^v��4v-`�h�U*��^i���������ސ��O�mS�7i���Zң2�!�ʀ�>�h6��XD����6��a=�m[�M��+��o�{��jq6�d�͓~���A�f�k���\Xi�3p�!����ͻ#lZ;w�nu_?y��4G��t��X���F��3�.=۟}���V�����������*��*S_%�N#�}�����b�椇�!b�:>X$�]n��BՋ]���O��j��Q�K��c�M�zt0�T�l$Ҧ5��u�[���6f���G���ܒg�yq~SOK����.J�����z�P�F�rS��G_Jtj���`�d�����=@�0��wcn�8����`�����������?�e������%��x�J�q}�����\�2���k�x5�����=zT	�vqfu:*e0���U�Ɛ�������$�V�msO���	'q��1�L�Y��q��98�σ�jD����.�\�>m]�N(�+JF� �ռ�|�&5�w�ɘ��$O $Xp�tA��]�9�y	�(}7��t���eqkC٬B�e��i;��;�f����O���'pDy���=�ڷz{{�U�8�1+�· |d�`Ct
;�OdV7��"D���\z��Q�"ufgq��8�;�sW����{%��;AxYz�n�D�hl'��lݠ|~vC�U�7*�N�]��a�>�	***�?;����^���8�C�|���q���� zm���D�pH�\ߣ���.u�Cv諎��`ȓ�ޏ!3�޸�C׼��@��^oe��W1��(�,�ruu���ه./{u�$rF�H�(��A�p�?2�ќa�xJ��$"D�X\��S�|E䩈�w��[���骯rA����}��T����	c���.g5'\���ާ��
MTO7���G��S{�1����<|�O�l����
Kޫ�k�%QWQ��?������z��6_���6Z��f����^Wm�.��ϸ$�0�W�W0�L��,����2��U��M7 ���0���ᶝ���(������#�~c���w#��N-��t�B)��>zl��ߦdV+|�	 �i,�f<8���16���in�4@�ر�o�x?�95���-�	�f��9F�o������r�����94�O����<Y��x���O���-2�s�DdeR�n~j3����3�gc������4�䬉z��I�Y�ٍ���+ �TU&�s�H�=�L�\k��C-�u	(ƻ�g׬vB֮�>����O^UrH����ga;����G!��5K�S���Ts\����ɘ�\:j|>{U	�����o��i���'�]7p�X����x1��}��DoFd6>�"�:��Ym��c��gli=�dA7zbSp�~b�@�?�[����#��A#l��;�c�)
����xP��7����������z�֟#��h��	�:8�zn�����D� зy1�{�ٯp#g,��G�ؙ5����>���,��������ɘq����5�\n���s?K�V����$�1�7�YѰ�	x��`Z���s`\~�J��
~��e��_<ϊ�P�pD��L��^���7:�}6�Ψ�ǐ2\koCX�G��3��q�)��<H�S�F�ӈ"�0�K���K�
g�F~�k��~AO��?�Ҍ��3	q�Ol�I�9&�E��zzf,�1ow������Tvz���|�Ljc_�ZQ�Uy��1B�y ��Ŗ����/�G�u�� -�<�ƿ���
�h�$hث�G�Z�p$��{F���f߂�۪���-��?�G �+[R4�ŀ�u�vw���
Cz��J����Z�|M�����6sA�����1��c8�~�ͬv�$��,�d�1�:�N��Ł�݉՟� ��Km�n�<���  �MA�jL(��:�kٯ3�`Q�}�$豵U�t0�rf!��g]��hn�]���e�^^�k0Fi��}�km|jf�23ҟ�R���FC=��3�V-C�+R"2@�� b�Y�����j��]}8n=����ZSX�k��[�� <�-^�������C�;�7��hGe������2t4vJ�{�l͂�-E�:%���ڬ�˙��� �܋�˔�}J��.����?u�do�������K�@9g�����c[
wuqY��Đ�y~}�������p��Q�;��g�%��w2+>�����ID����&m�?��\q������\2�?�e?����ask�����7}�q|���wà��N��C�l��683����C�cf��R;�p��~�
%ج��+*b*�Иd&[���{�p������|ļ��`�TYc�}����/[veuM���`?��K��s�7�﷏�.8��ӳ!"ݣ�C�ZV�Ǔ�R5P�߯�C��׎��rvn���}9�.��xJ�ec��
�֔�ŀ�]�n��P
��ql�Ū�� /w#^%6)h߅���fm�;+�,�� 1c죌ǻ�Cٯ�A&����g?����@��6_��v�7��vt.���k�y-���L$���%	Z�;�4�/=�(=���^�j:S�I\phX�}%���%��5��r�~��� PK   6��X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   6��X$�8�l  �  /   images/aa130aff-16e6-4627-9689-819d55b5861f.png�YUL
��Xq-EY܊����K���a�RtY�_����;��kq}����M2s�9�L2�3�/Z��X�XHHH��Jr�h��[0��Ÿxl���d������?�m����p���d��e�j�����e������ي���&�D�	�F_YN����3�z����k����Ԏ����(�Gǳ��R��7���c�JMNf������a�\w��{�I���kD�b�K@�)u+h��,?I9=̚;�����[�(6-�r�d��CGG�%��+��1A������G �����B���	�A�eF,M��Lo���k�=�8%_<�3��5���K4�AlaA��~��V����6�~nU���٤�:Ƌ]��d*
����W��CMy(%.KL�)�U~3"`��&���Y�t t�I� �Be���qkP��r�<f|0$L(��-+_�a�� m���$�J&�a���%���}$?�}}����4��ۏ��˜
|<gX��m�/���&�f27��+F�lȏf�{L�4d
�"��)"eN��_���`��N� �W��ܥ��d
ڵ��Ϳ:��-�^���X*�^�☈"G��oւ��^���i2���n	�ii��}I� ��M�L_�n
k|��g�^�D���Fg�Y�U��'�Ԥ��������$k_{���A��G�1�F\���uGLvaf��<V��W��f^���2=Wt���\C<�m&�	@�Z�O���g4��͆R����թ�#�7�Ȇ�A&��f�vf5
�"����0��hż_�z�@o*���I�3Mu�l#�c
���H�Z�I�C3n���6���ﴪ�	�,�@_�7���E_��~��ܫ�[&�N4�X��������'I��^��D��;�d C�uI'��;�����L��ږ��!�@7�<�^�����	�ʉ��!Zv�pt6�L(�QbG���Y��XHZ�e�<Z�L�$��K�V�jN]��{��i[E3<ӿ����R¼�`�ӡs@^��pv�Z�#�A��4d!~�D��޳%�{����i)�*7�CՐ��\,��{�_{A���>�Mu]hm�w�bD!�$_`�12Ő�Y�D	�,��&���W;��uo��oX���N��������c����`j������{���c�sH8�0'ޠ<C�ȲL�Q�ۗy�ߡ`��#��Q� ��y��IX��L�J�{�X3�̓0�1�|'��f�9�CC�U{�'T�K�c0�W�&O�BMJ�7&�꠰l�j��������X.7��k���leY#zu9`�4;��w�}U�@�l�`V�[�Zl|D`�eJm�c嶚��lnQ|l��;�l-��|�8�Z�-b�P˪W3��OIƭq�:��KS��d�iؤ�)��)hDסQ����UU��e�K��iKR��@�^9���� ���7G��*�p6�����Ir����1�q3��	
�Fl�I�=m�h	� }9!��m�W�:�1�jC�����w�(��b�������l7��2�~xJ�֛}���F\��w.5��ߔ�h)UV|il��;��cL�{K��ty��{ �``���C��p�w�kz�����I��g�'y�h=;�@�D�{:j^.�m⅊��|Ǚ9����;R�ȍ�� 3����xw\���CTl�y�,u�v�e����Y�(Tc4@X�l?��%:��v�M�(��� 8�TZ6�[��_��Rz�#�E)��i�{�5��.�X�uj}\m�w��~&�e/���H�8���Q�/���H�R��5���_�5�q��i�V��;���~�++�9Q����9=�CK�;G�T�N��㥲b�=;�p��>�3���W��.1���E�����|��Kv4/�t��XTJ��6�u{��%Ǻҟ.���G@���:� ��y%��
��E�N7(�� 2�-���]�H���Z�  O3�*韭�<m\�����t�pz�#�����Ց��Um���C�nĮ�$�e����uesM�����?����pc"a�4u�hi� L���(|�ϯI�L� f'�E"��*٩��ծ� 9�-]�]�������S�;iSKn`Uȏ�=����R��8�b�96K�A�E8�կD�h�⢛ns�/4��b�#5���6�R^&h`�j�y�9w�T��ێ�Gy�x˞�iz
z箹�c�*�_�9��Rg��U]���,.V�m
g�H ��rK[}����цQ�I��X�H�����rZ�y~ 
�6M��
򗢧���A7��!ܡ1�@��I�ĩ`!�j}���%h�	Hm=M��ğ2�2���I	��F��[�!�Myv�LE)v��� 3���>�xj�+�Ҹ��_��a^�h�$�ՖL����q�Rf�.��� ~D��O(h7G#�<qF�[)�������k�mFG7fL�o��k�1ջK����r�W��o���2Q	-��k�z�Phiѕ��"0����u��{���blRxk\�SK�.wFM=gx�)���;��(DCR���=���}���ST�P؜f���M��9M��X��Jlָ�.�1Bf�b�^�����g���H��(�_��_���	�F�(�P��}�y�&(�$՜D�Կ!u�y����e��a��,2�R;���ٯ��=����"3[	���6�rm�E?\L#vO0Q�3g��ˁ��m93X��GS�=]��F7/�=6��z�|�y��0�7�#�����7�}m���4t��`���H�袟���P�N�ɖ��{[���4xʨaO�K3\�qd`��R��sL$����;QE�I��G)o�LQ�uz+v׺,��L��X����%�\��p34p��Ѩ5 �j��Z��g�<6�^ܘ��岓d$^I�@//�!R}�V2qPN��H��b5~�q�@ ��>Jɒ��3��?9��yb�Yř��s���1]%���Pf���&O��O�X�����S���cܹlb��Ya��@E>��7X>�J,#�В��s�*.i�JeyL�P��N���	�@׾q��/"�M�))��u�:�����T؃ZV&���b��(��h5�]�+��9��0�Y`/��|�~�<�����d+�_?{����@�U��bꎘ�״$�P�`oP��R`]���;1�9<P���Ιd��`��rCF"���\ջ�(d>�M%DiJ+(63�Cb|"&��x�xL2%ѼZ����CV(�(�aW`��m��R�E�o�j�SX�r$�h�cz@�S��.������/���kW��z��[���z�K[�tK�f(��z�ôڛ�I�����r��,�*$��;$�|�q���zw���ǜMh =J�"2�Ƥ7���"Q6�˪]p̻�Aզ�s��:�C����w�5�hxa8B�L��n{�?���(�͸nu�$��Lt�z-=
>�EO��M� =�=�pΆ�0٠��Q��e�Q����_����h9>�Q�?O$W�d��/?-��uh�4���)(v�Uh��CJ���/Y+���<�!�Uw�~]PP�����Qǟ:�Ǟu��o0��|j�sv�%�U�d16͉-���Ze��Z�PR�_Y���7�������}���؆X����Q�������)6�	��N*.)>�.�G{��3�L^�u��p)��ÔA�Q��yM����Vp,}(Ll�xh�����---l�PT�ruru�ޥ2c:��n.1�N�\�4�M��3�ť�N,��f�e�����5i�@�Aɭ�-YQ�S���fƎz�
�*w�ÌO�ƪ�����'�J�/���#�%��.���U/��G�+;�ET|VP8�FBM����k�WY"���>ފ�]Rl2�T'�w���QK~���O���҃��b�15fBv���tA��g�q�<QӳRolև̅����A�D�.`7����B���*��R��$�ka]|o[d��J�=Q7�FbnO��I7#b�F���3�|�T�#1��D:��/MV�u��Be������u8T��'�&*�c��/C��̊�|b���,5|%���l�W�d�_���V�{������)���y��4C�dZ s���NX9�[T�W�⍪��ѵ� �"*SPÅ+W!��q#���[Z?��Vl���{�w���	�h�i6�XJ�/��I�\#�)짎��~��x����@�'^�u�! "F}���P�����@f�kM���������`mO��3���((��MƠ5g������본��N��_�b�mjВ��W�O�٩�7W�}I�.N���وa�lF���ʔG���N�$so��]�S�ee���=~뤶��@��N�z�5��:�s���ĕ����R���5֣o���laӗ0���>��^q�������3��2��R�7�$�;;M,ˈ����B�������`��W�p\4�\�qH��� `����1�T)!ؒ�Ak�J��b]��%{���DW$����~ս��F`(��ÑuCg��F�(�+g}}��'��- A��x���6����n���#<�]��a�������{�c��J�,�5�p��qp#��R�ZX�S�/.t�Zr�]A��a�N�(6���_km�mR�c$�<Qq��)~�+���f�Z*pk��Z�f�͞Ff�/eꝻ!Z�@�`ḋ,����?)�*��(�<E"�3/���"���"��o�{�RX�N��/�a��ZU���xm��iX21�:1}�,aS缈M�rwg�xM�u��k�Ѯ��e�k��V���S�Y2�֯�Tw������o���];��nf�/��ŧ�A��\��W�o�@��sފ�H�#��3��m��{"�E�Ӛ�G_�U�]��K�i�,�E���6��tl��$N�J�%9��{�P#6��䓏�#��.�^YSx��WBI���7m��O99.UϹ~!�t������	�[z~� SX]�"{��#���7��4w�M��z���$�o�,lM��u�D�Q���=429~� �����AŚ��Zo�Fc|��a>Bz��
?�.j}�"�F�4�'OdZ-�QB����j�IF���{$��dֵ~�l�EV&y�˩ XXy��DJ��c��_(}��s�T��Ҕ��[��D����Mfod��%������Y��cZ\���$�1�\�Tgp�ڊ��-��I��*p8�C��k��Sm6\�������<� qN�&,&L��0���=��M*�+Nol�X�V�ډ���b΂��z�o�����ӭ�������YĶ��U$��H��)�5�:eW���Z���<��c&j�0�b�m�վ�s���X�O�0!R+"����U%���a��b)�[����z5g��x�$����Ke�����d�@HN����c�܂ח��):__8�$���8�+�Y����JG�짽�4�E�^y��5p\���h��VU٥���h�븏����|��^����ЉO�I5'�V�t=`�},R*G���8Z�]��Bg�X8�F!�E�����t���2;ę����+ݘ�V��L�Cc}����)[�-�� .KfwG���<8^h@`!;��6ͮΒ��z�Z�%݆W�Z>;�[��#���0�%�o~���<;z5D�)a-��X߼}��U����[��̸��W>[��
���D&yY��~�}���cx�3��Ey�1�VC����wv�Ӝ�)1���Ⱦ��L=���V}8�LRo��N� <���5���w��x�4����O�߆��Hc���]H�Z	Qi�{�������ɳG�լٲJ�����̸�V4�$E�2�z�5�|�R�$5R�a�qL�qe��"V������X��	�y_6�IG�41��n����@l"�oz�i�v�ɤ��KlP�*$La��B��g4��i��/��<�:�\]/����d�!`7��k��J�AVf�����Pmܠm�g\|����"݇�P�B�?� �jdԇ�-�#u=
n��m9/.��\����\�]��g5<�����y4�#F��C!;I�@&0S#��T}���wd�@C��{�K�H1��7��,���M/�K>���-N<�6��"�wqN�5���s)��G�q*%���9L�Q��0�wk��w���x>0.A$���-�?�˙6/�PDH���>��2�P����Eiap�13.�U�Yz�C�)|�s�VkV����#(V�ʹK7�������ߗ3S��n��?�p���gҏ8��Bقo�'j���BbZ�%��M;#w�"�⮣c5~���/��IseIu�/�}�m14ƷS��b�#�<��k"Vj�͇�[���V�o묆I��?DoA	�Sv��&��������d�~����6��v��h��=�X�?mΜ��k{�����6�c���W�L}c�w�.�S�~�Y�s�_ٴF�u��;��8���g�����QT�0�ap2�;Z�1''����>���˵X�D�%!�$�ʽc��V�/&^+lB��IJ�(��y;����+<���V�ܮ����z���Evu:��2����=���!�K�[�xWK
�il�����qn��>I���-��UI�rub�j�=Qut9�{̝�#� Y���r��q}�V����� q�n��6f������O������e�� �b����`���g��8t��A�ש�x)n%�W�7'��C]$�3�������M�s���-|��f��9��A4K�l��@F���D�����,��ߜA��[/"*����%�="5=�He;�^	1#F�,"�e���Zo�^?TV����_��z�^ЦE>@�
>�$�RtF��1~vu>'��s��K��Wk�pϚq���A?\7�~ϟ�_�G!
����&h4�[���

d�.����g+�񿩧z�N �C+�ޛoxt��mS�j�����;�'���kpڜ�L�]��)V3�� ���R"�@(����l��t�O�;���;�
Yͣ>*'�a^9&۫]�g�7p�v��W�&�C����C�ޮ�����lloP�H�l���(�����X����}�`���cZ��S���h݋�e�9Am3�P�<(�L��ho�|�h.Ϲ�о'C���F�"�ʉ苃��7�Jpk�xsJ�3I�U�X��V�D���6 �OfQ)R�R������r�l�i��Q�u�)��-�a�5���D{j�b���5{f����컈@����㠸.;����}l���p~�;(�:�6���,�y��{?%�9민
�8=*��I�)is��c{�{�#diۥ��,��lhq���W�!��a s��[q������%�U�?J(e(�T�sZ�%�����>��RnӺ��j�ܿPs�>��l��n�wEl1�u��O�!D�	B��Z���bC�~�3Px0{�#�PR�_�L^��,����A�ǁG�	�?S�א+}�PK   6��X���7z  �  /   images/be8de2bb-09ef-440a-a2d8-19619bf9d0dd.pnge�uP����iv	Y:X%D$���e���T�[@���f)Ii�R)ARZ:�����>����s�g�{��3��+Z]U���PA���֨=�A��U83�t�7�@C���o�����B=������r����p�A����|���ae�j���n�u(J��FK� ����>�&j� ��"�>ݽ���vЦ;������p%̑���a�Է���Z��R�P�Źy����S�3�g��'iĞ�j�8�Z�%�Ww�G~ڝ�ջ��\1��pY�ӭ�Ǜ����L�>�����֣�I�'99y���������_�_�"�m�g[#�w�G��,���o\��%�*��&����o�i�7L/�f��;��`�Ҳ���>r�92��{�H$�s�٣���<??����QИ���?��)�G��5���>����7��II8 �_��ia���0-��;���>������r9�ﵗ� v��eE�|R���k?�-?=�l�o<�Cj�A��Ӳ	~�e�t��w�´������K(�
�\���.?a�D	�:����'@7ݬ���� ߽�����}aG��o�d5�J0�#�I�� GD��i��p!�X�x�l��G��@j>lF{�����O���`�'1�		��`kQ��k�n�+�߲֕VR���@H&����ѩ�_Ĵ��� w����[Tx���F�s*�m�E����N�*�]cX|�<���"�P\��҂G����ؕO�i
�=I�Ҩ�8��#J�h�6:N/-��ڇ�-N� 	o��Y� �����O�E��{�
�/���L�kp@�wy	d�Dލ�V�����M�O�ru�Ñ���7�M*�P&�i�$g�P����ơMؒ�?J�x�]�'6J-M��%	т���bq��6K*e'竏*��ӰM�%����[��w2��S��፮E�@y7�J`:��;��Є�>�L�Jq��1x��J�
�O��[y�mN�P���].�H�ԋ���k7�ܢF�G�u��`�e�Q����<$��v��a]A>4�6t��J�`���&���7k���sJ�=%Nm��	�烥��+g����\e�tC}ە�nsߗ�բxy9�WW+�IfQ����ȳ�ID����)t-�=	�(Ke�z��+O/L8��0LDQ6�P6�(�T8��C`�)��ڔ|Ox���˧!Y��u��`���8���[�}��f�/�\��S���8�\�����^���B���İ���B7[�2k�L�t/Ũg_1��ǃ����p�ҌI[�A\����&I��ϸ�G�������4�ihI�	CX8`�<!�����3���xnՎ}m�}��Hui�!�6��ޟ�^��D)��_�]��� ɴJ�+Ţ�ۅiiC��
_�$���b���BF�GHā3�%���㘂>�{:���,?�f=�i���$Ga��m�Lx B��Ha���8���݇�ǣ�4_�(U�&���fY-2F�'"�A�^Ui鱋�lB�!具�"ZX)��חI���r�6�9y�@�nj��Y�L��KvQ���� 0c�'�[����ǘ��1�ߔXb� �ٙ'�x�˓�q�
�b�������Hά0�A�8�.���nc,��|qrZ�ޖ�����+Gٽ$]�6&]��L�u/,d7P�����O��4��rtQ(�U7���[PX���Қ����t�����cp3�
͵\Q���l�;�n"�;����p��y��!�;����Zt�f��>jg��ƾ=��O/�^���TY�� `#o���t�L���QD�����-��}��B�M��es���wh�Ϻʩh3im_�6Yb���lc�y����]�0�Cw���0"�M�2n;��85{���Mݱ7��uҵ`|%A�z!}���
i�VT"�X��e>'�}�	ռӲ�H±���l���b}�?W��qɄ�������E�W�M |��L"�!�2WW������tcPh���wDpo�F�P6nh�����[���a}��I#{^��X�p��ŌN[��j��*Q�==�%<2���;,r��$���7��_�k��ƚР��
ݪ�Fs�S�}[�|W�eG��������~�n�"Do6�K��u%����a�E8��F�D|��2��C���5�^��q������<O���ƹA��s��(��4��(gp���9U�0���޳���TTFHQZj���z�`�k����	Y^�-e%�ˠ���܀Û�����Dq{y#�r��G9�2I��"�Ke@;WҪB�y���hF�z��TL7�&�ȨD5�2K�> �Z
8�OfQyw�'�!�2�q��-o=lq�E�O+�˭�X��'n{�^YOI���v����y_�V��o��)�\q3?Kf���^��T��l��]�Tӯ5�Z˗~q4��#���W�`�����Z�������ed8>%�Y)-�	� ���'�;���$g���)0�Fǔ;`K���l (���y���S��O��߼�>��r�sQ��l6<njڛt�!
��<[mg���s Bude��g����1�\��"�}�&��2?���'K'"��/$b��o�2v��j��{���y�0j��C��3ngZ�;�6�`�ݜ$;��TJ1>�jll���8�6a,|��F�]�ٹ���۟�;��V�Vqנ/���õynG�jo�M�+�ݧ§��~��'��I�4�^O�����H��/Qδ�!����jz3�����͙�b=6$���nE�{��k'v��s���)���`�E���i�g2#�C�=Jj�MO2�����z�֡�?h��F��8��y�&l~�R\-h3U/�q�������������K�h��|�����X�I��r2F�54H'��O#(�Tf��*?�و�����}��"%�����ۯr]�C{����T3����0��6��{�Z�h=��~cdr�go��Įj����g���3���f�z�g�[&�GՉQ[. �WNn�wU�o.�#P����$t���!� {z�ѐ��s��L&�_pgk��d3��[��]p��d�*q'����wUN#(U������~o�0�����g���J8�rC�@g��%֤K}a�( �؍�Vy��%V���(d�ru޻�����q;��]�J�W�a�~�&��L3r�a׫n(*��l"9����t'0�@�fE������t>���Uen7���i�3-�7Hw�Ol��;�����L&L*�qLoFJ��?dǰ����H[5^(����+1$=�\���e�9�L�^�^b.s"vY2�j�|�Z��6y�n�J�E��j�i"�����kd�|��"�a� ���J�����B�F���4d뢦@;�7T�K���a��x�Ǆl��!y
6���	�,QjK�f�3�	~�X�)X����K�[�h掲�4O Ϸ���V]KV2���<�/�pn� ^N���. )��r�׀AᏉ�<�C\Á�}���Z���G��ˀ޺����v�N�"�W�ȅ�؊���ʎp�&{������*p��BZ�!(���������(�[�S�13�i��"P�%$w�Dd2c��[�k�Dώ�ǚ���ux������`�����͇����Q��
�4�T�f�k-���;��)����^��Mc�*���ggҊ�գ�n� SE6N��n~�iP�/�[q���ʮ-v܅y�R�ˮ���뷖�����efx��C�N���ɽM�O�gq.?���ֱ`�ь�ăz��'bSrԍ����to�7#���F�a/�C`�e��V����^ZF
]~p���6q��$r�`��$`�@��N���y��%5���#�P����ڬ^�C�q� 0��)S��2p5=�����d2���g�Wb�>C�&���]�Fހ~�Hl�G�����!~�UU�F4��魕��]��#�rNWN��r�~E�Ԁ���x����ݛ�:SUB�+�*Al:��}���P\����1���C�uRO\�K��X�}����6�be�~�ܶ�_�x��8y�iL�L�\�^�܎B1s�,<o'��=��$<����(�a�8[�B�Qe��c�3��4Y�Ҧ/�u��	T<?�N��F���r��|~��6X5A�H�;��5mЄ�Y�޴�m�A�eU�9���VtU���G��{ؼmX��6���tT��J�m����e�x�4�Mۇ},�n2�H�.E�����ʥ��Ftv?���f�[��H��.Z�;9j�Z�����t��~����e��V�K�*ߎAq�D��,�1TP�Fm��c�
��z-��]����6�eX�������l{�U�=N�u\:�M���]M]�T6�c���(��:<&���!�w<�q�� �F�s
�6� �`��|ѐ�
�����L�����qbЏ��1w��;�i ��7:Ќ�_�?����B�{���F-�`d1AcQ�o,�b��Y 5�d�{��A�l�������;��_�U		'��=;f��?�U�	��5�|��������oWtp�F����t' Yi���g��4�L\C�[�r$�	n��4�F��μ4�;h��ޫS��W[4�[��u�jX�>uW����G��ٯ&���ۚҗ�X9�?�Ur�<�6�O��'�[�F��_^Vj�)7c�1�z�s��0�����oRrNq��t���f�8_Q��2H��q$?��AY�j9��p�_�{�U�6����-��DMn�u�z&?�ϸӮ�dk`��Ķ9��_Ā��iA�5��yv����ꋶ���M娖~,.��^�gį?����J�a���%Yz��v��#K˸�������*C���}�Hx�ټr:/����\��,^�A�y��n��k����>^7�t�L��'�
D':�ϒ����/oٺN7�]����}�j,)Ѿ�R��ɲ�<�2"���	Ym=�pXG��-IgN����KT�lukL�>����L=�Z�zAC�D�F��VZ�q*��'��������Zd���6��7��g�M:�7^X��Z���h�!��Ŭ메"X������x�9A�6�	��O��4
e3���h��zDxg?)��Y_�(D���,49�jN$��˚ůE�C�	g�Qe��f�{z�0j�Nr�̡�9�s?j@Ǳ��Ml�����C\�n��{��9�ۡBھ� 
��t}����|��Bl�t$�#7��57���~����Q� Ll�d��ͽ8#� �1S�_?�1p���������-�JZ���]N1�Wߗ��9�pP���@�?Z����3�U������H]�'��(5�F�kx�<�@���qbM�qZ���(�����|������i�A�n�<&D�V��̒���x%0��=���u���y���h�����kӶ���K��v����yMc�t��8ZvR���֪z�~ń'��rb^����w��{�$� }�i�R��*|eciN��<`��Z-����0�U_��e�3���K�s�֠W�]�M�%�hh��)����fO�3M1��b)��?�]��l''�M����sTBKӨ�4�׵�j��
�����9y��ऻ�����j~�iF�T�M���k��>�����3Wo�`A:�FH����X��p�>��
�/�ii̮����g�DU<�&&͚��L������,(=��+F�:�E�,�0]޾8֗+�_<b�|}���u����X�^j���cL��5�Qb������Yytl��k�ǨLM=��?�/wĉIX=#t��qxG"t#��*ΟY�]�t��7�1��_#җl�U�S��q����d��g&t�znn\��{,!�)B��q�P�P��p��K��M�	��޶��C��μ{B�ZHR���x�X�OS^T������9�x�sS��$����R��ǹB̬��F�1>z|65l����M��h7,��>�ٱ��2�۴QBb�(9Rz����ϲ��>���e�������%�z�8(s�IS&�/hDu5��o��r�%(Z�
���;�ρ@�S]��,R������ڬJ��@!�_��4ƒch���%ѓ^R�6ihJV��٨��{��`��t�\FΥ�E_��+�le��_�o�E'��V�MmE���B��������5FClwh���&�3�;J�K��X���HM|ląv��K��D4y��-��������[�V�~���<Ź�@����7�:I�j����H*N�W%J9�P��O}Q�Kj?�Ո6l���>݉�g�����r	^�S;�~;"���Տ��z�n�f�2�����XBDF�ڦ&Fީ�����>{��58�QkH�';�:�1-Clx��t��i��)W�X
( i�ޙ��2�Ow��9?�׏��0�-G6bdN(�����7�Y�~�{l�vz�������mg5\�#{�����0�N���3������\F��7�H��rTD3S�~s2������:`�8�ER�,�;��[���mtܻ�ݫY�!��w2CS�ܻ!�>vK`���Uf,�&��xH��,9]��c�b�h��R{���8o��K��z���
�y+I�Z.t�Ӽ��:q~W�Pzh�Ֆa�Bɻ���
����+k�]�|Ȫ��H�U���5{O��ǔ|�I�͡��^	��Y+N2W���"�S���V-$�{)O~�����g�;5��d/"@���J��W��txnh�EU���Z��.YL��<G�3�
'��!::�'�J��؉/�Z��F��-1�͸��>�������M0BV��ہ#ׂו!����|���D�Ko�<�EY�4J��mZ�5ԓ�n*��R_�|LMܫ�\�Xr���(�bx� �(��SK��t�2�|�x��]5�Ey�KI�i��c�A���K������������=�	����h�U͡����*�f��� PK   6��X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   6��X�GDU7� �� /   images/d628d844-ce42-4e82-be63-f5fdfa438334.png�wTTٷ.Z6ݢ�@w+���6�d$g[D$�䌒s��
[��,Qr�PD%I���"�Ud(
��Cy��w����1�p��[ٵ֚�ߜ+P��T�~��+�����1q����u�,��oT���g�����{��%���Ώ�����3-6������k8Y�#��Z �H$������gn'W�D��5�O����5���?�9t	��T�;N���h?ڏ���h?ڏ���h?ڏ���h?���-`�9����t졚֏���h?ڏ���h?ڏ���h?ڏ���h�W�����w�>�d��c̯��nq�������\<W�^�)�����WvK��[���<���N��s����vK`_���jv�z�n�����[�o��p3�=E;G�oZU�y#3�{��4�.�����o$��0�5"���x���ȏ���h?ڏ���h?���Vh^���a=)n�$�pX޿���g�\�+S�(�6��](Ӏ	�N㱒�w�'ӪJ�����K!�:Z#�|��fXN�Ĳ�_���F�cv�n�|�؝v��T��m�"���2��/�r�f
y���f��XH����S�V����z��y!�R/󘭮3���g��o �3����Z]fk�>�)IN���;���n>����9�}M_iX�X
$��D���������+��\����4�ͩ<Ƨ4Ƨ���)?�Բ��W�`T�SY�V��o�j���$������eObՕ\���Ն'�k���_��_*K���5�\��ubK$��G�0 ƓT�g �\���	��i5O<�yfMQ
%��ޛȻ�T�����ښDq���F�{L�ڈVav��>Z�f���Ԑ���dC��^��?���~����~Z=Ͽ��%.�
�d��m�%����_�)��$��e�9��LM��#����s>s����4Ҩ�S�n{��)���i)���;�z�ֈv(�]sh!:�v��|7����e?�o��O{�'�T$!Ћ3b�V@^n;^Z��K^~_jҤO{j�/kM���u�<+F�K��)��{yY�T�������^0��,Sy�/x1j�N`!�X��6'C�c!sB�]����E=	��CMf��]:퍹����jؤ�gq��c<�����Q��.V�Ϣ�e�C�J�TʌquoA���Gs�������3�9-C�퍽.��>�ٞc�}���E�'���q���~gJ��^,�)G�M�O=&KyA,�$k5�呕�������.���5�9�Ӹ�?��6 �jf�����5��� ���˔��l�2[���	x���r����!-y�79'�f(K��Ȉ�cl�� ������]�R�?�g��EW�󝲯�l�]��B���(�	Q[�%h�yM^X����/{�kF���Xy�ZӤ|*p�W=~�
k����N��s�?*�K�.?.�KGi���>4��w��r
�C�'�8ܖb��W���Ȝ"iIS������)�3���/�c�^ֿ�����?�;�,XF
��ߋ�T�:e�b2`ȴÏE�n�m����.	��Y�Cj-S}�22���k��ͬp��@8A�(^Z߼-�H����$u�l�rg�a��,�:2#�'6���ϭ|��j��^�>��=�G�O)�*Yf��mڎ���FT���)CM��4Ly�'���>G�=:Iqc�0N����M��9{��I~Sf'�߅�=�WV=�,�9��Bed�H��Hbל���KN�%{_/����bo<��K�X��0n��U�����}��8f��
h{�춡+1#�f����Q��!Y� �!�~9/{
V2�����qK
n���X8<�#(c�!(O��m�G
� x<׎���������W���Q��T;4�����3���~6HB���ۄo�.��BF8�l�0��ܹ��G�d]y,��Q�Gx��8�oVSR(>'��q}�%�"�L	�5�#8���R��z�����`K���t��AygP�����A��yB�#'M�S�=q<�5�t�N#=�� ��|t�t����tS��r�w,�h"��J��\��.��mW48,:r����[C�":�ڠw��ˤ����Z?�������DIx�j�s�Fk)ec)��!#�矂f�e����ؐ :�7�&��l3� ����	D՜����~��x��`������BM��	�A��]���&�R��l�Q�ZD��G̅�,V�
�5Ͷ�"�&�����F�-�4���Țm�&����6�\z�Y��8������WF�y�×�����٤3J@��g5��ne��ʧZ@B'=֙��(��QÆ=���u"��ƫe��0����t�pt�����(�wL2Z�B@#��}�ݯ���HЫQ���Y�k�g%��Ǹ_l,�p<~�q���s�U��	�����<��k��9�J�7a��%�ԉo���y,��v�*&�?d���\͗�o�~�b?g�}d�џ�S���X����M��p"���������4�d��<k�z*q�A[���R1]��h��Ē��F.afG�ec/@Q=�mt�|&�caK��q;������_;�?#m�u��I���*_�U�+�ىPo�<�?��9�
�:Z%Y�G���6��^Kt�) +���/Ol��S"N[ɤ�~h�d=�n���;#ЮB��C���I�����	�|�`/Na�z=�w�s}�#q:F�����d-�F�\�b�����r;�kM���d�� b�B�q�
�hd���ȡ��k��5��]�Z|�F(>� x��+獩���"��꽡ͲZ�Y��:�m �w���-��|J���:xH����rC�p�b�@#���+�2sy����Ȧ2�וAu�"[�y�Hm'��};���� 7����z6-�L�ג�E�V�5Z��,S�-���9���JEF/,�hx�4��6�T�cޜ���z~��j���I�oGNoS���{h�͛q�v�~BW�O���	N5��≡p���Qdw@�?��	��¡�9Ц�PL�u���9{�F�v��k�z����iw8��_�P���5�@Pkհ�����_���(j�����Ԙ��5e�5�np�`�':2{���`�/���fج�NwbĂ�Ưz�����drQzDʆ�����u�B�N�z�d�{�T��9݄jy/��v��F�	��G	`cS�����-Czk�<38jOM!n����RKg8�wZH�J8{>�a�r=��^���ί�i��g�}���k1��Ff(�D�=�kQ����>�;�m�x��k����|\q_���
�*fy��ZDK����R���*i睬��I-n{+�y*� �X5�Z�Ū�����|��Q��34ఠ��0���T��[��P���Y(��Rr&�6�!��m�J��kV�])�f��t���?��n?/���`��I �f�����X.U��_�蹤�O/���ʻ�����X��¢ʚ܊��E���*�ApZ���<&�
��9����ƻ_:��6��P=�"���OD|�}�8&3���VT�x}�>a�}�ԑW_�7� }��]�kP��T�,�_�$��J��)���>��Ĕ�����f �r�:N�������gf�m,�&�h$�y���AM�% [!t��b�hz���$�9U\S�Hַ��7�©�����!���m��fs�%���}�n��:�ǖ𲃃߾���Yd�X��݃�A����I5�c��Қ� ���`�y-�vG_�F�^m����q`���U#&#�>0�λkK�����tGP��_�@�'"`�w�	2�d`�NBv���e�����,%�q��+A]��X8��tҗ�a0�r�	FU'����� ���K��%N�A���B;��w8Y\��u���ZB	CBl�Bi�T}��4����!n��!GF> $J�v9�v
����?Ɨ��qF��j���_��CwW�zl6���ԛr�@ 'L'gY���?3��O ��`��*��r�� ��W6%;�VzO��~�+/oP���1z$�}B��'ȵ��%Xc���@τZ��;Y�Di���ݮ[^�cQ�SYv�/ݰu��.�V"P�V�!�Vˆ��h����]�MM?�%uN(e�.�,��l���[�4q�+�oON/�] 0�޹�f�
�x�V������i�ow�Tp�Y�#@N��Ax)���.6�!Њ�;X󶁷�}i6��XeH��#�D)�}��V��k�Sⅅ�D���v�U)��$�����P�c��_A��d�,FQ��E�5����&�K:��s�g�&Q�}�da�aay& a/� YO���F@�$�I�&�#c�Cy��&�Z�u�x�Ƹh��~����/�1+2���%�Gx�%_z
ՉJ���`*
}���G��n3�,��$}�~�n�n�Y��ӵƷ�G<&M[XU�S`�:)c��H��#�_����fd��|ڝڷ�'2�;�\,�jP��� ����0����:�
/�dGGZ�!�q!׋�&)G[q�9)R;<��SNb�ኇ�1����o��>E�&!�֡��ޱTc��F�I������s6�s��R�<9Ҽ�Gc���	����bU4�/F���1��V�.��~m]p?��������� ��"�,sٗ��F;�QBF�=a^Z ����P!S�T-'�f�8����A1݇�$*�Vf06C��M�ƒ�do�A��R��W���fc�3�> �m�wq&�\��e�N<p |n Ӏ ��3�:�f����r�"ڽH�0n�;�$
@�
v;�Ku�H���j=���-��_�ç���F%˞�7\�PQ5-���!�n�"��?�?*�ҷ�-������P����_����Tu�,��?E*}�5��V�.�p�#v9"���3�%��	�R
���'@�Dޙ�����M7�T�o�X)�Z`�����ܞ) ��HX���)�/� ���i��jʨTt����f��e�?@���~�هIo'�)l�(��..y�1�yǔb���_�]w��{{�[]�t��4����N���K&bȓ���� ��]_!n�u@7��s��eW
 �V�E�ǆ��_�;�ӏ�����HR�H�c��/u%���!�b�)����=������:�F���YO��9~:��� !{L�$��O����Wڨ�F��v5��'p�a��;�m�!�
z^�"PH�G}������k5�U�FU��[�%�8�H����o�2��8�uиa-��f�.*	u����X��j�]q��7С�!�,���η�!�=}�����2����qK5���6���;�;���d�: ǝ����:��/s�en��u]���S1�F�Ě�b0p�Y�R�e
�/H)! 6�L�%L#�ч[d81p�[��~i��@��h��)�x�M�~��}t��V/J��eS���lޔ�p�����DT��"�Y��$��2dٗ�l��׎��LT�e�g�H�_�����a큏��I��$�?Y�� �Q"����HȍJ�F���QɅ������,$��򇕑��Ɇ�Z��kl�>��HUyW�Ң/�:4��&L<�������6&:���<&�<B�;����P���Ϩ�B_li��E�K:*t6��e��n����8�f8�b��Í=��j���4�^$]�����	;�=oL� rp?��L]q��L�<
��;k�j�=�p6dk��{�2�gS1�����>Nr��7�#��ןBR&��Rm��tc`<���Ȕ/4C�U��"���X&J�O������o�U��;���]��%�;�r�!�YC�/�U�H#n�'�+W�k�j	�'lO���1)(㽸���<cFZ#�!���lϔ:�F���cJ�PqE�:✯@B�man��R�+�"�E���9�/�0؆��� [��l��w��R×����:������ ف�s���m� ؑ�����0�H Y�h�!k	���*w|Qу���K҉��f�t�﮿�@)8��q��+�r��j	���Ie��)�ۡ�LX>up�ك�xC���q����k:��bZ'��p�Ƌ�A �D_������y��k;�|�f�h.�9��6.�s���zl�p{�1�GR-���v��h�H4����ґ&��o� �����2��0u��6�rHI�Q[og�*6,N�Q 4�$K�x�&���;(_@-T��ӎ�Oy�{9��h
� �)s'�NR}M�jiCxC���G�R$�pe7�G�e`ŉ��B	{z:�q@T?,�58�;�U K�R�$fd��Ԯ&4�ǉ����p��#�f���(ӷthA���[���-W��p����j�� ���0b���+��B<9�D e�;MMdL|Z�໽(��-h�x�H��^�j��2���>#4/��u>�����R�/����=N''%D<A��pM^���z �`n����o���ete��4����DRX_�v6�é�IJ�����ƳnC�_�#Ƞ��M�7
Oړ�Z�f%�3����5��nӰ��rk����,Ɩ<+4�? s_�C����%����+�y��P� �޿~�V��S�N}�̩
Y��S�RQBNÅQ�>�����h���g�d���D�Z�� ��X��U�D9 E�j���r���	��!fA	)�������Zqwh�n3�ސe�jû����G�ztp�CLA���r;�ѳ���6��<P$�9h�L��[��/��o���fj�� ��ɻ��#q$j���2Dv�Ԕ�
�O��<]��}�s����օ��T�����mD+�lha
���n�S-iUuzOjK:$��B�B����>��8��%���PZUI��绛i7����i��\+|����1���^����q�<����������x�͛J��
�������+u���p�� �V�T�SBCu�x4U�/U���|��5aF�xw_��;��=Q���f!T<����%o@fU�+��~ ,�2������w�L|����{��0����/Y͚pjܫ6�+��c�&���=2<&Z� ��� >8Х�sa��3~��7}�pV��&��m�g�^�-KG鐱������,(W�d�f����n�������$!�SF!��hNڽb��t�72М��p<��[L�����ca;O'�S]�Z��$Zi���:ӇϽmv�M�}�,/`�|̠.�@�n�U~�����h���[.�}���>��M;!��ܪ�sQ�i�����P�?u���Ӿ�̴��������:vE���z���͌UU5���GN���l���;`"���Hٟ6���űY8:�wA���]'�Z�����o*S�i@�vv�ȎԬ�_��G����D-��)���R.�3���e�����X���l�Ӗ4�\QWʁKK�Gv��)sR����Г�)�{Y�K�~ӊaշ��=�n�σajJ]���k-��&Q��H6ĩ�ݴ���5<N�lA��OH�6��kJ�]c�W�@��x����H�f�'R�ǖ�9�!:�0�o�MN���$���``�@�D�ξ
���T�y�ogϝ,x�q�d�$Md��w[M� cL�NO�g�(:�唛���L��13��,_	���Z�-l�����@2\��p�&�+�&�2u�J_��u6��9\۽�u�|]Ľ'6�H-�E��&�mf��y�:� ���z�,g�se� {��
�.f\؎MD&{��߇٬	�M�X�Q=U�Ho���.Ąͻ�
	���s;�nB�?a�L��5�����4����/>�K�7��}�������a]T�_�+���5�)qB#�w=��?�-~3�k������5iz�*Бj��fVc~�bI�X\����2��&a_�Eq�er�d�Gͮ����=j��r{+�'��<��{�n�з:��7�6T��i�9��L��Y(GTw��8���E�i�q��i�'2kKLV����������+sP=5�M����.�M�Oږ�yKQxJ�P*b��(��qR�׈�2�Oe��pe�CM�r��fx�֨��N���@������2�7u�%o������=`���$6���"��}� JHFҲ0}j��6L��(�n��S�`u���8���
�M���@�(�4.G u�
��)�+b���b��j^���I��)�X���.��i�FD7]Fڝ�X'n�2�!�d��/���	�N��d��XD�3��l!׾�ۻ�m��Ś � "^�9�5N«���C�xVט�y� ��o¤##�b��Ò��8|�À�!��m��rq�vW��g�{�
j��=Ӱ��uk�@o����[k v�r����5���9h��>�4�����z�#>�S�8�3|��G2Q���A)y
&�!Α���T~���o�aC�\MH,�]��Oߡ88y�������`uL��bAw���sY�����9���ԝ�2���od��^~�"j˖��9`m�(7c���t�/��:��tbl�/eU\,��N��Z}��y�R$z���ג��Pi^��U�禤I)w#�˽�!�[�Vh	�Z%=^i;�D6�d����e�Wr��VQ�R=?���]�M^kr�='�	�<븡�Jcm�r;P?ry@�	/bB�vo)����"!�0�t8�=l��gaS���Y`���NLT6�n9�j��Cb5��@VU���zA�� �){�J��u� �Մ�'�
�%��p��@I���1{�*x�J��6�Jɟ��>�c�o*w���S 	Ӥ���B�K�Y<�|�fN�D�����0��Ǉ����۫w`sXFy�tӈ��)��5ښ�
XJ��*zۖ�%}%���{��UB#��m�[�s�O����)��keDڴ���B����ה{E%g`h�oڀ?x� Q�^C��ȿ4&���0�k3�ةxB��&+mN���DCs�+!��G�մT|X����.�ڞL>8*F��|�?#���q��G!2m�����,_T���b��SjtaP`������^�ʛ��R
7����h�
�%~��0:�g�Z���ӷ�l� �/�W���&�i�d�;��Z�֣��V'�G�7��_Ϟy	�L����\��w�ӱK}#�)��5@C�#�3;ycT�o�����_�:ё71��#F���+
���B>�tON�������M-m8�Jk�=7f�g�`?���TX�Og�d:O�ߥ
\3��\�6V�+�z��{irn��"��ʞc��R��v�y����`r����K�4p��yQ��Z���Qȳ�C����HXL���t­�~��T��J�~�i�l�t�h�N�r�jo�����`z���
�k�Ȧ�B�QN���-5��*N���7��Ve���*&k�	iᰲ�2�Rg�`�M�U5yr&�����j��a<\վ��o���p��z_�������s䶻�@Q�]��x��c2r�~+Z*��k�Hl�2�]0ji�4S���{v4+b��Ն�W_QF*v�Eބ�� �����Ya�O�%���w�7���u�cW����:�������j��]J>�,?�D�j�2]�5��l�J��qx�qz�@���C��=���H�>��x�~��Po �:��Vf�4Y���gz�ܦ^�kK�Jy�!l�d:� ���A �x`gUMRYPhp������t���A�nTN�~1�lb���n����I��� ���h"�â1�n-� ƽ��d�-ݡg{�N/+�JV��)���U�kgz��a	k=ˣ���gV��!�M��	G��݃�D���� '�/��$Jx�b�T!�gL��mz�qÑ;�u{���h�����  ��	CgH��_�5V�O��-H�U���0ғ��TDU��8� m;�L�U)#�|��rimRî�S��)gn~��81�t
'm�XV(6VV�OF9H�n��=�M���v�����;'�i�oV�Y{�2�rx������`c�pG�����^��K��+�e:[;n�T@����n�T��	���I�&3��9�QeGQ�j+7�Y��<�u�fR�Ǧ����d�	�J+�W��j��S��	���z4T:�3����ۇ3 19t=�쫩X��Q�@�f,���2�f�7�KB�"|7
�H0���@��w%z�w+ZԷ'��]=Aw��Y�0+�m}n������JK&Hi3(hEd�Hp�>��#���Ѧ��"-�F��5��!��
g�y&��A�:;���|��������UE��g~�g^l{����9�����Y�b6��f-��c-K��=?:��Z(ͦ`�kLs��/���1�q�/p�6�;��8��=��ڃ�!4����Y�_,2ȵ�a��`��]�A��>e���lj{S��a��CG�����@uv�������@ɷ�D�e".�Hp!���K����NI�;~�pg�A�jA8�a�28Y@�ޅ[�"����rF/C�:��nPg�)*'���ΛVY�+ʄ2L9M�����<�9a�3���Ϊ�uʧ�
Jѧ>}�g)�:i���v9j�F�'�w�^��;��q�(N3��Uk���
����-Җv^�f�0`Mw�
W�#�jBY8}U0.�΅�p�9�#�xJG2R{gx�i^o�Mp�s�Ag�Уw�cq0h�{�f��5Nn��A�,�:2�C�&v��n*H�I�o�����qU�,O Sc�d��6��&O�#@�.��䨝�~�������Jܛ
��k31f�!��%B�y�����TVQ�8Dǝ����y'3ݪ�OP���1��ĬQ�ݼ8&��Ғo�蠂����}-.�_}����yk�؍b�bI5l�bG�̙p����t��?��%,a��6Jo���yN�8��t����� E��1:�Y1�'��������L*�J����δ͝��>&y�.��mF��o%�����O��)�]�I��G��?�3��iuI�Rk�(���+ez�W�AN��\U9e���0]V��e�ɚhS��W ��̊�S�|����3�{�\�����L�r�Ɍ��i��>l�qwY��Z��u��S�A�%i� 4r�9h��|Qnn�I!��v4�2��q�����Jp}-�0��K����%�}�y�Y6�+�p�6��@�3�3�K�n([V�`��)�
�t$L�U�+��#��sܧ\���fm���7�e+?{O��&~�Rö?�E��?��8��3�?���5���|4Um���/�6��o����fR}e�[_lc+��f�C|�����Q�>���]��+�'��Χ��DH��� i�h�@�����#$�I��o �j�����Fm�4�)��x��f$���h��=�;e��z��Y�U������ �v�B�-Y"/���b�a`�{=��8���"���_K�=�,W�`�AKq�Zez���\�t��r�>2w&����XT�S�~��^%\��CWC:�u�Pj��3؎*�O�c҉Li�"����PY�h�hق��zF)x?s덷,qʳc���A^p���2P/e��{�C{���"!{@�a��H	���6�-8b�Hx���u�#��yՍ>K��՚%�?�_y�;Ej���W��7�������e�]�8S�0���
&{�Q���[�4͚��L�*N鎘��]?/�\�)��|(�%��$H[�U�ꀷ��~�u�NE����X7 �h�w�+>1*����DE�	�#*��p�WU��U�*i�#g}�"Ȃ��ދ&+���l��\چ�g�~��'Xg���7�{��j��K<;I >|�KR�n��K�6�M���t;㙘������>�1�@{�-a��r����Zc3����!�+lT{�N�$RǤmѢ�ddD��y�'�'������Dl?2�e�H�s��'0{< W���8��d���[��.˪���;t�zˤ8�s����t*K��]v�d���&dbd*��4��坠?^%�U��Ԉ��M�'j�Aoܫ���
R�Do�sA�!�&*�?Q�ؙ	ތb���b�t!c.��jx{:w�<)�k�uj�k�&�����R2S���7�i*�N6K�ٙ�Mn�����X��s� $��%z��}�D�S�Y0j3�%.��8o������Y�
��R�zn�@��:�J�"��'˴�!����"���D��
��ӽјyv�G�z���i7J��	�A��)(|���X�Avw������b� ��n������+h�P����J�L�J�N:Y�c$*�)W����0Y��I.;]�&��k_��p��5:=�>��1�tv!�:���T���C�s�����=��@��"y�����x}�
r�� 0@�[�_�1����$x���b
��SKF��*!-�G'�: B ���9|m�L�f��'��6���S@e��Хjƾv��|��A�/�L�n@�M������
�#IYC����11Xs�ob�=#�}̫��PJb#|��m0�g8�m�����&�¥�:�T��`���T����̀AiGB�?φ�O��D� ���۸�7cS���F�\J�}��*�"`ę�;��K����������x��������� ?5��-��$�;�O�Ƴ9y`��'��cv�17�)�Z�ջ��8'���F��2Ż\�\�q����:"�z_�������&��/������J�M�'�o�ċ �ԡi������(��������L<NFa���{M�j��X1��<�1;�Y%.9���=U���j��`ڮ���} !�j��v$��p���:h�%l�nY�]@���C������cx^ӏ܂��W%U��)�6��䭦���e��2�$[�K�s�Q�����c����A3�{��l�C��%=9ЬV�@�>YW���a<�-!��� 
�He1��犹��&j=M�:�=�P����Yo^� #{"��q����~�o���Ō�~V_����X�j���tl�/�&)Î��&{q��Ϋ�fo�E�a���t�t,tJ�ae���v`��\"�X4�N�w1��C���cR1-�.24�^��ȕ�kr�������˂փ�Z���?�d����
�����-��}����L��.�i��5n�X����`�{��CU\vW0f%)E͛�e �z�=�̙���=M�[;OF*>q�<���a�2��3
�g{^8Ѱ�v�6�� �d+�~��a�	�����8�!J�����W ���v�Z����NJ��-�h���o��z0[�n�A����Y�hYYh�. ϵ�>����2N�̯�1���zoj!B��3�2^\?2�%��ש����.�r���6f]>�~[�+�XBh`��t*��X�W���O�J�A��-���\!1Y�!aM/�'��ύ���V6�����H��`CO�v�)N��]�9úڙF������<�� pz��p�&����Ƃ����%�/Z�:B�5�W�Ғ,Y2�cg&1��9f���=�O�`��5�I��W˒Wy�_`���s��w�(�F[�~)��8(��;:a��������G�Q*R�t@IlY�8�n(���Ơ����6E����ʑ��]����n�����W0�
h�H�P던ٮ/�+t����]D��;%�.�Z��D�������jt�6^��;T�[���2�׶[����5k�kUŨ>*�b'�)t���چ����ai��n��(�k	��q 	�X��!����W7_�ܜa��<6"3"���3��F7��T�Tn�Ak��;�	�'Vv��/pXs�w�ȫr��p�:m��k�A	+��9���.,L�ݲ������\�[��v2Lq�ם2�>cG[z��)�mo�p�2�Oz�������k��exr�aW���)�*`�/�<�{��HLL��i�V� x75���3u������0P�4+U�L�-��<��o�?3�L`��������S����%`��	����.����	�ap���r:�u��8n22��LĢ����� �3���
6�"z����7������:'=ԟ,�ήDȽ=�N�@5=��s�>�Y��'�I{�,�f6+t�+[o�<�)��Ѣ��ݥj��@v��d��W�~O!�ݧʖvb��V_�Zo�<D��� ��V	��z�\���
J�lS
=�?Q3��Ь!�B&G���)oGv#M��ahhz�]5b��l�֋Y�2W\r���|�����"�/c0㣟��I-�����5���O�݆��?#�!�I4Cqdx�}f�j�z�O%L�j]���"	Sǝ���!��'��U�&�J���4���pqU<w��2�{�2
k 6\	��[��̪��BKॹ�;��,�s��r�]n���T�����`{����j����b�*�ʡ=�l��&I��5�%���Á����-i��|��^H�`(�=:v���]�`'Tw�$?�@�oL?[3��49����D�C�dU��yō?�Xn����l�9I�u�6�Җ.O8�$���e)	�\�@�o� \w{���f�I
>�����X��OA��gm�X�͍9Ζ�3��:\f�.fgҿ�����`B=C1\�&��ݏV�$���"E��"�o� 8�"�����tA��#if�>[# ���׆��}_�:��NM��8c�'��L��I���u�:��?�cu��)��T?�� ����Nd{��t��;e�������	1�t�s��+�-��������������78�,⼕�Jzb"���6ۏ�۪�
������k���=-\۴]����B䏷ѭ����l#+��@�P`&�䴇X�z�?x�4�_���V��h�&�s���}�X@ʚ/SKTw�{���Z��D�L�Jh���է-ȃ[&��:L�Nˑ�O|���-���4
4�&#��n��Z\}N�Z@�y�u�3S�����'�;=CQ�(˻��ҥZ�/���m�[�b��k��������8b�G����;r�Wj�x�ᗝ�͡_̢pxR8����̤2j[9�dC1�vۡ�mt��sj�4����O��3��&ӱbko��y<�H0x7x�K6=首B�\{˶��d�q+����V
�`(�o��~�
l�U3���l`[�O�;�������>L�,�7n����{���%�{6�C���VJHD��?��W�v��R���3�N�:ĭ1W��y脏'\9��t��y]�ZR��h6T���]�z��dqg{`0CX�_��X�eĤ�Fh|yU�T,{+��`��ٿ���F�^��f�����{��A��C�q��;P@{	��SMF6��m�jD.�r,Q��O��}��4S�b	bXHhx�?�aB��9�N�:C�/|��/��4��d0�{_�'��K���fO�r�V����gF�s0{�'��Yl.^��ؚ�,; q�~%74Y��F�*�����:5.-Ѥ�s����s|��?ް��
0�z��\�~��bJ��G��ՠ{���*��v�j�/����o�~'-��]�1�/�����1���N����5�9`ִ�Q���~R�ڃbؖ�%/�o��� ���h�0B#ɇ֞F�ݎe�ޒ˿8�<�*u�8(�/;!li(@�����4�s��w�R�1�*AϰgNE�}��	<��
es�y��=�q�_�8�ݗ901�.$i�7"}V��0��2�x��BKY��g�_������Ƃ�n�{7v<���?!Ď�f��D�B��7ό�S�@2�/�Y=��m�C�G�7_��3f�|�şu|��~�s��<sW\v�&��(�$�����7�ߥm��)���%%F��)�쵌{)�-�~'�{���=��r{�=]��"�G�D�c=������3!�cv���ps�*���93?-�'o��a)��r����{����p�86[˵��[b�6�q����#��t���Ӽ����2�Y��'�i����Ҿ1�t6
HM]����5O��en�Sld��b+k18B5YA7�k!���,:*��W�ĥ��ڽ垈D���!6��>�)�|��}U�B7�k�=v�.A�A��lC��p��� ��&���N͘��%�^������-�A����[�3�_��+�h��D}�ʽ
����w�ఊ��]�F�Q��"��Ho�j�8M���wv9۰�ٝ" �ꂢq�aҡ�~�RN�ߥ��*F���O��P���`|�y4
�����E9)��[i��A2$���ۗ[�Uyp���Qb�̬[`c�/�d��YOƑts{�l�7��y���nH4>�Ҽs��%�+.F�R��x���nJ!���܆���&XSB����Z���vO�M5@�rkȦc�f)��ft+D���������aŮ��x��C�Ql��ˬ���l��M���,��"z�~*r�@
S-�(�Xt$.O�������_T
v�
�E]0ʪ��b�sN��ދ�p��`4)�r������Rv�y'N������HVzV�؆�C�o�C���9�{��=?$����` �����ۅiξ���F��l��J�jn3@��o��4���G]Ɨ��D�:J���J��9�Wߒ�?�p�&Ӭ���w��HT�Qi%W]��8���$ߦxY��S`��$��k@�8:����ހZm�i�t�+F0�eD�!���+�ަbBXj?n��.vrՎtF/��u<t�6��0�Ap�%����sզ�����]G�oU[���������%h]F�]1���~��I7鲺eOR1d�ψqP*�٥�4���w"����aV�Y���n6�~�{ĥ��_$oQ$�o��,f
g�jX��3#+м���p���>P��#Dv�[ᕈ�7/�$dً�OR(�/T�	���=�:h��Y�\�d�\�1"G����G�������.�#$5G���e��ܕ��A38�䵙����Z�5��xQ�k��1S�
�I��xf{0m��M�bW���
�����5�̽�w�����BUn��%��ԭ�����uߠ�;��	���U�o1�^��+O,"���QW���6���~5��}Y�������2������D�{L㾃IS�����?O?�9>.����_}������OJ�=��u?^��i�3��Hl�q���ɻ�L�
��qו�O��FR_q���Xt{�Z�\�?���<DL5�u�3�YP���s�x�o��L}���ʽ�<D@���S�r����ؿ�f`�;J�e�i�
�?e/n�.$t�Vbq5Y^�g�C�շ��O:X&���з��}����"6I�=��T6�w�C�KD@�ҷ�RYN�(%&[.�>L�����uB4KD#1H��?�*x2h�5��7�5KH"�g�ʅ���*l�|�\�
��)L}�"����%[Z��I��`���ց�����o�;Ța�_d��h�x�6��N�o��1g��:;���of��'�`! l/R�ĒA���9y�ĒK������Bĉ�s���hd��Ա��B@(R�s���T�N	�
.t �c@'2���;�fd�oE ��Dc���'L�D)p�X��]�����O�N��Ab Ckyo<h�,C�ݦ#�
ñ$���
'�T��X�&}aCOQQ�I����6��~~{8�T�[i��D>'9Y�J��[���wgμ�j�����v�,V�t�f��5O��]�L�hA�������tZ��j%�����-�U�Ċ�O?�X���q�/�����{�]j9X�p!+zg�Ej&��2���d���u����-[��m��z<%,�6݋[ԬY�W�*F��I�z������Csu,J�ɑ��yW���^�gBz�n�� �D���{��!������ATT	�R:��Hw7H7C�
R�Jw]J���!9t�{����>�~Թ��}�^{�}�=7~�	�j�oC3f�i81 �H���W�#��cV���7��?�!v�ŧ�=J4N�VOh{���	��DjT�N���Rd���b$���J�J=�XC��I��=�G�X�d�r�:EL�& ��$)����,�*A�k��6�����/M��]4� �yuǀ��#�5Rt�CiE�Ѓ�U�6��i>-?o�m:�!tU_���A�=N�5��(�ME��!Uh�A6�]�[���J���ƹC�X����^5��Ĳ��-� z�3�z?��T��8�c-w��E�����ط*�&S��R�������S:��_ ���ƴ��+���؂'pU�`D��p@��hקּ[!{�p��"tu��f�MT�-��D�9������t顸�o�����Nge�飯�e���zrݡq��A4/�1ʣ0���p5��t���G�8��Dȶ���L��u���X�8�ẽ���%j{q� :���l&�.l,�<5ta{���$˟�{����5@l�ʪ����{��hX���Jo#"XA}kh6l�L��q5�tn���s����*%���{0�u �����k^+2����M�R"w�*/M�$��:����ޓ������[���*���=��!��� �"�Nʴ;AJ�2cǋ�LG���웗�xth�AOmΙ�o�K@�e�k��IZ9�-	��|�)t���H�I���.�����θ�\�{I�8�J_��5J�����ا�g��G�w���I|�5:M���)��Aj�ġX�z�3�c�[��+nƲ�ܩ�k��R�N��a�r�HrS ś-%t����.c�
w]�`�G���Ӡ�b�i����&��0��a��\�U��� �V��K5�3 Oj<���=���Ņ��tm�g�܀�ȣz�����s�_�,����*"����d�/X3!#�<-׼&���m��� 88����VMJ5,վ�`�����em�����;���z�~;�z�$k݉��;/!�����]T��TI��%����&�\�ڢ�����SCbp�(v@�l����:o�͟�V�I�u����]л�����!����?�a�<�'��p����ޱv{g�⵵2dM!f��� ks��6�t^��^U�)�����4bg���>���&���w�ݣ-(�q�m�:`C'�<�t1t�9�-O���M�I�AX!VS-,��r^q��RzwO��x����1
Թ
�ߕ��%�T���/�<R�?|�H����o�q!2������9P��T:YQ^;s���/�Ї^���Hrx�ݿ��.� 9$P�
gp���T�]�P��H
�,6f�����i�UH��he:͂tBhe�3NCZ�I3(-�:24���!:�QD��M"�xԥ�^/.�6�LT�&8)Q�+6y����J��o/ �'��>g�jd*d;���y��*[�h�(�z`n6�{[�P�J�'�ښ�V�|��!��������(e��eҶ(���r����o�Az��q�+�]w�Gu/��x@���T��B��5(�g4����ᦦt�׼������s�4( ��U�W�P���(���F��f(���?Z����b�"y�\ƨ��E���Q���Jd�V����k��]��� �?��>bX����le;fM���̥�G:�O��.��rH`b�s���%t����5W���r#�_N6?2U�`G=*�8���,����B�H}�Lb�.�Π��~i�O,7h�`)��o�o���^��8$H{�q��a�4.���;,QҾY�vl��ŻJj��J>M���^��2+R��c�>�B�E�0SA�2V�~�΄q[�@�l�TJ�k�����*o΂w��4i��
w��9�.�!Ζ���ܵ�	?Giv��o�&��F��Z@7�	��&8�l�c\T�+�?��������L�"�X������23:����m3J^���6��\�s�%X�Q��޸/v����ib�;n� RHu'uµ�r~�r���Ͼ�-�}�L⌲K�{Wm��0�/�ڃ�V�j�(�o��w�=}��=�o���e�Vn){�Jx� H�=�8"J]��՚'�v-�����l��r7%ݎ��5���P���W�����6�����2Z<��	��w���L�?�+�	��_=r��L=���@[-m�Ŗ���Mo���_�S��Oᕭ�A�Qu�t����K���z�>�ѵ��y_o�bR62�������%�xj.��Q���a���eB�민�]�����^�kMoן�/���-�9��:�侮=7<�J&��OY�0��-���/���-�@(��m�B�ᣝj1�fk�=������s^LT�o�`�H�A!���)��	����Wo�+����)����jI_���tR�7�Y:=h �`���U�=���'�6/]�-�Sd_���r�#���H��<5b��W��R����C�^&�~-�p1f�o��������?�`0g��?�<�����$�Q���6��؞X9I�������2_��	��0�dD֘�]���7�D�%X�/5�5ܧ
��ރ�;��D,�K�w]d��c�-0��9Gm��H���݋�ͭ3D�-z��f�����xy���_�*��E��80Z�V�e�ܑ��1�-�6C��'�����J��?��\3�f/:���%D�^\>ޏ��#���)�����?��`�e�Ѹge~�ypt�3�6G�1k��

ñ}9�o��4ǰ�hP����`��p�$	K�S���*���ڛ����b�~>��(\u�!²�QMB%��<L���:H�>��h�~�(:��N��-���M�x� I��|�g����.�j�,,�w��;��ɾ@��]�=�#ԥ\�y�v4+�b7ER�˲jaڲ�Z>�y[�Y�n������]Mu�U;H��$��P�#T+�O�˱Y��}ek�(��%R�O~��k6vڛ\�z���Q� ��>�f0�Mݟֿ��ٔ���M+��d��W�~>�����~s��'q�'��V� ]��;�9y6��7Θ��6�9�.	~Lr���Atu�_����P_����� v�.<�E�Ǵ��������ƕ5��4�]4�y�����+�ɖv�QUɣb�g����H�qh�!mãp�;8�|捔W�RK�#�^����; ,��<����n1���-�����6&�z���۬X!�Ş6�>��A�r,���x��7h߾�{��{;QKA~��}R�Ӣ�}}�7d�~B��� }���ϣg��:A7�{p�������������w�y����M��
�ʎG�꺣��!�Ş6$��6�5:�DV�	���5����^��O��R4�_r���m �x���]� �����y�������:n��	U��j͒ʖn�'�͖�)0}Fq�U�I��\jBf���#]B�G?�t�63���{ϼMg$Ĳ?"�ر�&V�# S">-`GX9�\���f+M��9�+�_� ��4p�PňPw�@�K��b�|�Z)�ƅ����a:��	rbӯY��ո����4(K��:�z&��u���ݟ�Y�J�iy�ۯ�Qc��;��#�XaH3��ł%��zu�(�{f�l���ˑ`�׍֚�`tٍ2 ��>Xߵ�_��@��׺�j����肥�<@� �t�&ߙ֒I���Uͤ@�]�μ�p����L�yy�D��f���I�e���c��R:e���4j�Wia��S��ԵV^o:�۳u5H�|�[�,��,���-s���Ȭ~���~�E	���
Td�MLcj����S�|���i�o�C��7����V���}���}��p�X����E"f��O��~��������e6xA(}�¶@Y������XI�/-?Շ�.?�f"~)(׿�V���8}\��PU�(E��eǠ5>�38<��I����
���[�5m�Oט�g]n�<6o8�oq����]t����%y��D�(J8�%�{],�X�u-%s�I��A�����2Y'�/74���C���(?��t��I&>���2-�ĩj��{E�{L���<o��菙WMx��{��e��S������=9ՂX̏X!K���Z�1��Fqa��ه%}�h�� )�=�7��d疏�*)�T�]\�GQ+j��cQ2l�>x9d��T/%܁��lձ�����o䷘�E������s���Y�(�ò��l��X|ak/^�)��B͍����an����!�Z�>h@��dw��F^#�+�~�����\�n����o��g�Gٺ�$'9��K0A��t�� ��ujVhPns��py[ӌv�9�p�<�W�:�3~�����C=^�ogk�"�� ��I�C�H��U�n�QA��j!t�H�Ǣ0=G��x�O��'<`����d��'"5(T�6���Kn�5�J4��t��^�7[������.���
P0�E�ﯤY�?.^����7O1��t�*���a/�1@�j�f�hԚx'�Fg����a �A�&�,�7�r��"9����?����I�tH���H�TX��d�w�M���G+���҇^n�ALbȶl�V=m!�;�AƢ������>{k�H��<(�e�߳��G���f�j���k�\�aU�xaؑ�j�$!��n�a�oĩ�|ޙ��7(/1P`�#�	^p䏄<��'�͉���ﴔ:�Y�>(Λ}�VXUc�JȎ���g5��m���>	u�;3�/������I�jf�xؐ�l�L�)��F+��O�x���y�|J+��%)�(���G��7��)�K4G�*��lͳ�p��g߆�ɛ	��w�x-76轷BTr4n[#��M����PF=�b�������@_����@}������iH�M6�d��U�P5cɓ1+# �J�:T��o����v�k�����oWwj��!TǊ%R�1K�m�{�񝻒~3e�]���Gc�~�k^)]70�~�d�Ԝ"\Q��u�3 P�+��k�o�/|p}�:ݝ�l8����ک7��a4�Ԑ#��_����`rOfN�;p;�A�R�觔	w�qt��ʽw���� ���ͣ�/M����	K�����V?{D���&	Pa�����W�஀l��`^��E��G՛]�Mp�!_v_E�Z�����_$Y�e�L,X���D�RT������Ь���2���O?��Q���^�:hɣ�RAGq�gq���[ET��Z*�a���O�g���� ��Ǫe�~��Meu#8�~�����f+Y\iH��m�,��d8H��:�D>b���X���UHQ���޻vX��QV� C���w}�xD�b�%�n<��DJ�PYd��0<�g�J��K�C�oA�����D�3n�C8�����x �|f�qE��SUr�% �N�{�1`V�W�]~�%@^�F7l8�IR;bV���l�v��~����wv�����6'�Jߎ��>�{��^܅�$E�7H��ͣ4L�C����1�&&/Z�������/�`^֭mC��;�t<~kH=B�۝���;�{k{ё��@{��*L0��'�uw�k��{����º}*<���4���p@ZhR[M�U	���L��	
e��j�����$����4ɜ���;��������*5f�煫b��ªx�G/MƊ?ho���0� w�;�_�&��Y��7�jP��Zm��e�D��,��G�Ga]���в��b,��y	�U���ü����%}l�I}MA���~0�=�	S[)L(�z9�wjc�6 ��}��'�*f��P5�.Rظ�dvM<~V�PiP~%!M_m�w�X1���|���W_��	��D�<{~hG\�#��m%�Pnm�!rl6���dƊ�ؓ�֞ow�zVYa�A���ث���D�V"���d�H�OGq�G�a-����F�Lڠǫ����r���]�����7H�*��f�w�F���+���"������n�W)Qm?�a�{Ǽ�B�֜�[w���),\��+��"vO��c#�Q�{�b��"����jl����;����������iI�9_G�X��K�Bgtt�ݡ�yYUGe,��|.,n��֢��
g����r�ܜr��r�^+eԓ���;�c��T=�.�dR.����zK箕���v���竄U	S�N��4������2m��S��N��׃��-x�=X���_ ��h��s��� Ds=�7E\k�d�9߭\���# u�le>�͕�ſv�*w̋Ö"V2�$l5��^�^�Sgl�[�s��N�h�R��tn3��h&?�����>��o=a�.�^��\�f��ż��ݨ���q����D�9��;c�F'�t��Fv�qa?.�+����j�D=���is�����UZw��n~�i�PxE��gz`��;nU3|y��$�����E����=����jʄ��t�k�|$X�e8�c%#�X�����Ht�G�ol�@դL�Q�
%*)C������Q����+�`�pKT/r�b�������bP����3�-���/ZO	�@-P�->i�Ns�Z(}
�?���zb��Ј����0rP�.V�ro���*��z(������+I�xJ^������>���0�[Y�^��=�����_3x�Di����������T��q!�|�J;�]dY~eg����)�i��QO������r%��?�N}��5�GJ!k�FƂ?�Mf8n�`H�j.>XB�����f;Q�� (K}s�YP���]�M�	`/����������w�>��O��'�����mz$�J6�G���k�C�Ϙ��cP����g ���N�^$W��QA�,u�f�����O(}G��&}����v���=?�|��Z�N�W�%�����{��2b O���bc���'Р74DN\4gk0��>����O�Z̭C �� �sd�jP�[�q�CAM�2-�S�9�k��������)�ּ	Z��Y��_�bg؆l������Щ��Ic�%����"�@I,�  ���.m�Ͻ�q�rlAG:M�N`�?#�R4G���CY7�৘���l����:n�0K� BW�^}��'�D���t��spR�0|l=tDXz��Ǳ.��c�>��.�Nl����=f;��v.|0����O��?,�=GM��z�x ����������[^�^f��Bd�)��巉�ER���#�w�.�m_�#sj�a�x����Ve�U��x�x]Ȟ�7�^eװoH��KC{�^�q��v�~��Br���5/���R��%��� �ǹ����W��������cn��}&F�2К�-lʴ�
LN�H,���g>�q��_�
.��oS��
�Ᾱ�ϙ�p��&d��I�^�Soh��Ɵh^LU%��by�:������*��`���j*IS��#-ٴ ��P�h�ʂ7�u�����ok r�i��σG�n?ol��nj���l�γ�/��H;?�U�G���?V.��g��|�j�_:��CҠ aњ#�#��9�
k\�eC_D{��d����,��ok�-��GG�zG^f�����w�1mPe,1L�tK��u��|764�MF���@��OGIe�Wj���3!�0�;�g���}å(m��A�7%���s-*���6~7���%~R�< =T�s�`F�sEgo��_�n����'�ִ�o>%�0�Y��tj,��A�~`зn�TFY\קQW1l�pz�l�4r�"]�/��a�\P�'c�A�fr�OPڂu�'H��.�5{oH�B7���������>���4���C%ƪ�a��@��=�����s�"!J��i*�D����3/�("��)��o`9EF%�m.�m!]`��H��웲[��VO�/P�,���~s��Q[��\��ocߴ������eHO��.|8dA��M���Mu5TG-�]�bmf��>8_Tr�C4c�
Y6.�4yz\�I�Z>~�g&��&�0�k�	�x��M������&'��ٙ(���_���� ;���L�;C�$��������aj荪K�	��m� �N{���O����7�ǣ����/�=���L�FP�J�����.A����R���]�B��j�g�+�#N�����O�fOp���xO�Y������OU�E3Y�!^^���k@���٬�5��}�Rme�\��{z�k�j�$7\��;D���Y~<Ll��{}k�X�p�U�DB�Pwh�ta�u���O�����²�����B3k�$���kȂ[3��`�m�� \`�-Q7HgA�diw{:�GMf`�W��GF�.���
�u%.�R�m	&��T�͠�������� <���[W]l��=8�s	�5<8qt@4U��Y���D���J�����������(��'�&�!BҍM��{��v���f�tb����e
� $}�NL���� �\�����Ypۜ�7�N��r��W@D�+�t$\�OI��;���E���
���	M���lA]�]�\�W����J��}B�p�L�П�>12�c�A���E�8�MT�2$�7(��o
��E��U=���J�$��Z����Q��t��}@���4�ɻ�+�_���6��I�����I��ųDa֒����<q���'�����{c�K��}2���ᡡx�t�M7d?��Y>��%��F�%G	h��kh�(�����T~�4�z��b��)h�_�ߒ�h�Я�q%�=���{���i{�FA�7�"������V�X�s�r/����$;�]��L���}��9�K����Sߋ�qr<�6�mB���ښ,����	��B��NA�������ѣ�|j�s12�]����v��Q�v�{��p�����A��O����������<��,
|720���X*Г�W����ݭ�%�)�����p���f�q/��}��~����9��I�2�е;�)n0)F0U�a�6�)�Ǿ��&�M�.z�lP��Ļ���e�gS O�!`���N\%c�i�+�������;խ_��b;�Z� �L.��\:�����:����ܰx�ӻ�����,#�V�gZ���l���6����c#)��	���`i>;�-\��Y]:%�Z���W9;�ڲAK`��먳Q�#t��9�&<����-�|G8���r��F��o�3bf-��Da�5B�E�K/<>��!���.�������
YG;��F�9Lo���U��X#\n7:"d�����N ���vOs;ȳn�)�w ��]�p��HԢ�p7H.YK���i�83�������H��[��a���5,G [�G�b���y�6[�3y�2�D9��\mU���3i�߮�&����(��w:����,}Vȇ��R��$�O���=̐&��8�NF�����em�-aչ�؅�
�(�*��������P)�+J<�;c#gb��3ЀZ\�G����:�4i���3)�vd��$ �]��'t9pC�X��8{f����~�hR��o~�zǪ'Dѥx��C򌧾�<�I	�0av9eӏ�M)�|ڦ	���޿Ia�����2B�Ρ�C�w�XW�b�����/���=8a�Z�zd�k]�|�_�^��>�|��/
;���F���"c{���^/0@��o����Y�1�1,
M��]�؁Ң�*��+/Ei��8e֬�%�P����ۓ�+���W��GQ���
�{,1���la�k�1K�,LrU�t0�8�����f�~\�Xb9��0���!��$��tM������3�T�Kj���f�o�,&Nm�=�Y;���5I�we~`��1�X�=�ڣ��B�MVK[Y��f�&��U�K��<�<[�ǜ���zK�"1u�s|�͏��,)��o�mt�/����C5��zU6��D]����Ok&��N�_�Ҟ�&�n�i6�71^y�σu{�X�Qh�_�	(6����l����=a�I�Ez=:�����%l�Iͨb)���,v)Ġ?�.ye��,�d�Ɠ��
��-��QoC6cr���(�,)2~t�7s�m�@��0�TڗO��$�z�0�Ӹ=a�˛ȧC0v�^C��	{�2�+.��*?`��+�m��.�E��歚C�����ֲrA\{#��7t�fLct�2�b�җa6d��{_	��ڛT��K3��?S7{�u7o�e�J�~��-��ß����B�\A^��;�E���R����m?�K:�Z�]YT�C�Q�vz��R�x�XjGœM ���n�O�$��u�oW����ĭrl.���/#�����Vo
��x�)�b�V���^���Д5�gN՗�p{pΈ^�F�%����s��Y���|]�建�0�k�+U��eEn�	&��˻.�HjfH]5U��~����^��+���8#�qq`�1v�Ҏ���C[�h�k��q��<q�����Z��,/�K���g~����5ɢ�c���-���bh��3�ԭ��XгK�=�G֞
�1��Z���h��yyy�L��O9����?�פ'$4�5���q|�i<J�亽+pL�9WCm�F)v-^)���`�`��?�^�ag�n���j&E���vvFEQ����M" ���=u,���x�4�ſ:W�ẘV
S�+����U>Z�-���cy<x0λv�y���9�k����xz�V�j'�VV���R�]��}X�à\
��n�a<�=_j��ܞNU��kˣ��Z6�*b����\�{D�p�\'��!��V���*�ESZG1�LP�c�y,��fh�R�AtB�j�t�ʃ.mo�{��Pc.���J��۞>'ӈ(�QV7���;��F�QU��y��-j���m�~PG�|�>n�kn*�e�#fz�4��LE-�(� ���V�/~��?R�(�Ms�K%����e�L��d`w��Z����/���ݗC���G�O�G��d	���j9դ*"�"~S�.���gv�p>��P%��r{Z=��"���l1��e��ֽ�;+�[��}u�ׇ�x̥�*�0lN}<Y�,�t��Lw�[Uəu�K�>�si۷Ծ�^�̻��#�UC
��9y>V�v���)W���B���e
A�q��H�6����?�Lds��"ڐ�v;Y?*��й�=�|y��U��(��Q����o󋨶�a���\6�IP&`R���5/���_�d���oyA�:^ʆn��Y������^�P����|Qji*+�ɟ���L ��L�Hy/K{?@�{��b��s�~E��f��lJ#�7��\��\
�t24�./����qR������m�E�F���-ѫ^��SOMwI�X�-�`щ��<�pW����LA����?��6 05;�1GU��P����
-L�ܾ����14{N��Sk]7,��s�=�;�1S�Of��WW12�˩�P��o���ƆEmJ�G�|�Aڃ�4T�X05���5�C	4k[p����C5�Ч�r��$8J8�~���H�����L����^���j�YܒO���(�]P6�H��=ef~�������"� ���/�^�����pU�'S��|�C��_X��ܷ�_�æά�$9x]�%���vv~.�y;f�f+<�zy�]xP��)�A��l�R�39�%�	:R��<��&-��alGQ���	��ߞ�W">Աh;L��`S�>Ĉ�w$0���j�#�Bѽo 7���Rr�q#�u�V4���ON��[#�PowS��5�������!}c���ӎ�C���iU��Y��HĆ�C}R��P�	7���7�ӕfɈ�l'P�L4��G�l�o���f��J����Q����K�����U��]g~������ψ���y^K���B�w�w)�s��q�k��M�ĩ�L|���{����κ{S?����ԥb�`����|�و	��Z��|t���;0�X󽱝5�?��P��m������4"�^M^�cc`.���=KN��r��W����O��3$e�i���L{��S�}�;����"���ꃮT~m��	uy%@�b�@��KG�'��#���N��m�'�/�b�$���E��5���y��^��i1\�8�)�$y���� ��IZ��/�Co�Y<���`�����6h���������;��q`����'�|����WH���itF�A}�2���F�M�}�Zhz�@H���v�Q#�\��T����ud��\�k&���*V+���.�<�G�n�x�Cb�;��t�6�P�kXW x=�e?V�@ނ�ꍪ���/H>m	���A�#�ݎذ'_����#��~@v�,0r)�}`w�ķ���S���ݼ�P`��f["��d@e>1R�P��h`��emeM�����,�}om�����T��%mE1�Gߔ�9Ʊ�v��ؚܑ�#pߔ '��V��m�l9?�Pk?Z�.D�R�_]���;�$o���h�4��-p��ޒ�V�m��΋�>�۾n�dgU����x��Sh�$�_��șZf3�R�:��C�5�x�	�k:���L1��kv�4���&���ֹ~k��HVz��\S�(���d���idY�e3e�1x�o�iʒ��վ�_H卌�͸�W�1�y�M��9k�$>m����i� �\��5Y��w�]d�e�I6���;0P�?c(�����zR�kӇ����"�r��FҶ��ʿ��a7�9V'�L�;a���?t���(������j����gPVف�W��q�$92�A�	� ��^8]Y=8&E�k�E0��I�p�}��!����RU`����7�����;G�5�L�U�P�k�.g��K�wK�o��8�, ͑�m������ ��Յ��J�#�X:��p� qVS�����s���2����h�H�O�N��ȯ��U�X�*�������>?��D�(҇����ǅ�1��D���pr�>��ŗ��*���mOA2��.Z�К�Cy�ޟEcB49X��(�Z�HZ�fZ�Ju��f���_6�6H�8��dǠ��ɮ�*�x��8�Ã�eo5Y��M�հ T����r,���8��J��AV���ʜ�H�.#m?$�%�~�4��)'�;H]�t'qCMF��a��*�L?�@���o���T�dʅX��a��S�Ĩ�8�}�����!���5��}�!%B��[D1Ι71���N^My�<��U�V����\�qTL�Ov��Z2��7�g��ݍ-��B~���%���R3���+Y�9??��fe<Es3mZ��'
�������6���C��������V�&��gf����Gm�Zd���4!�b�B�]i_�N8���\��$6���� �1�j&���v���Rr+ܠt%�X�W���ͥ�x�zꕱ�,���T[,����d��9�����¸��w���ކ?�y@1N�7��B��J?$L�Nu��F�H*���LA0��a�j(Q+Q��o��� �}���0ƹ�����)���1����Q���k�2l��	KҮ�̄�Ȼ������u�n�����H��z�0�'�f}@�
rA&��"��*�.b=��./�Ŷ*�V��k˵WPa�l�C
�]�KU')U*A��x�+�6�Y�mI���w�]�L�2B�Deި\#�3ɔn��j��~��ӕ����{v~��҆&}`��ּQ)O�������#T1��C
arn���E���}CP�m=�3)>�h��+��{2bZ�R��C����a��Ո:o�m1[�f����M&*%JT�TRn�~t�쾢��be�Wjf�0��.��y;�'n�w��O�E�F|��ld&�Zʘ��m��R6Z	Ǯv0_���Ft׆g	�u�O�%��3*�|�u�B��<P3F/`��;�'��ƾc����e��8e�F�Íd��~e��T���r�Ԙ����{MN%�T��Q�O���F��v��U�D�>��76�8�����$俯Ҁ����Ŀߣu*�I�R���2V�����aa$�l�_W�?Y~�kޤ<�tW�6K&��yHo��;uv�SQ,Ϫ�Ang�X��3�RC��R�G˰�� �ogK,fm���^L��3�J�E�\��0,�w�'
[(�?؛�*3�Zd~ �l\��r�Rvŋ�Rb��×w�w2��P� ,�!�
c�X��/���D�zc��b���ؙ/��YH�47�
Oɘƨt��^�W!\`����hG��x�Y@"w�M6W��k����e_G8��)-��1L/��c���@Pf�<��V�.E���>�p1?��u��gzr�c"HR3ܬ���`\G�IcX`�X�I�Ӱ Tef���<<́%����cc��I���07�p�>�W=d���\����o;
MO��	��^�m+����Ll�������A1 ��B'�9��.K��6����3[�*�%��`��~,L�������K�vVh�IO����hF���W��0BX�f�f��gM�p�R!�e|������`"�n�Fж�wZB5»o}�u{]v��I�Q�7�����2���S���D�s��Gv����ɠB��
��f��H���1Q����WܩN;ʁ�(�\���t]��#�Up0��դ�dp��R��5h_\/S1L#H�{�e�)`�ݣ����#Vu��%R:��F5�>!۾��˩��A]@���Ͱٝ]f��tFｈ�5 �ZI�S�`��>�`�E��U���$�jbK��[����Z;�Dd궷��� 1�P�A��pW6�~o�>�W����XzNd�O���H�r'4���������e��+�FH��@���RDNC����Y�Y�i;���5�*�O�d���9ޕ�g
�Y���e<11&4.��7v�7�j�7��*=�5TAkR�[�8E5���'Lob�����n��v�!��� ��c�lyE�@�l���K	��@���G])7E��>|�e9��4t�n�b�=�=a���U�d=R����Q��qR�U�n'jo�R��C��V��^��*�X3��u�Fu��Ah����#t���T�J>�Q,5{�!�½�*8�%?t��)jlG�J�#K{Gь�]f'�{�����x�I����ޤN.˟��UJ�BĢ��h�~v�Э�a��d3&"
�tP���h�L�u&@xn_tW�>���ȅ�d�;�����K�\�f���Je��ߟ.��)FP�X����'L��4_��Dy@�q�C-��w@]�r�r��2�A��Y" k�;�Xز5���;�⤟�5v�?bQֺN�V���Fz5;/�~���γ0�Y$$����s����׷=����o	$���KZA��5+��p�0MZ��N�;_M�\~w����V㋨K���3��,�vț���9�X �V+yOҬE:�e&?���Σ3ϡ⭹+9U2�U����"| �~t���y(Vl9}��W��b�W�;�\�c�ò��U,�ml�B��"ݺ�AD�j+��1�9������g��+��3�c���l����w�2�/%g��^nG"��!N|{[1om�������A9w+ʒ�T��]���ȯr�9I��~��Xh�{$rtjE5�	�? ��J�H���ņz�$w�g���v�*���L"D�V��;����L��(�M�8�l%�&��W]�A�W�Ki��wK�4e��L�ȿok�V���o�Û�eǙq�q�ȝ�ޕE���N}2�` 5Y�M������}kw��gj�a/��,n"����{����2Kl�͝9��fړ�e�$ᆽ�`;.���iIe)�Y��8��գ ��8X�SK���d�!�@���������~�m�0�@��/���d��y?�8iFF��S\/��}�I��^�ު�"&�OA�&�7�O�*	ZdV��eA��p�6l�^��B��I]��O���O�.}�\O)ܭ�t:��Ô<�-or��K�t�A�Ǌ!��Sj�,�G蔓�����KF=f�顈�oy|?��qx�*[�i&+��(*z�T�u�u�T��O��9hF,�T��g>�۟���]:���V�b�h����_����&��떁3�zPᏍG�	��r�wV�1��Օw�4�:Zs�s�v��H�F�B���?{I�,�����m��]:�O=�����l�����r �񘓧#��'ϝ�cz^��f8�P8^]%*\�~U�Z��]	/���ʯ�cPΆB�U~<���"��\�2���<���+��+�K�bm���=��\x,�3���3-�V�V0��6��A�����n�D����j~;x`%gс�?�HA�d�M�/�o��$��*rEW������c��:C]�5=T����3���3��C�Å#�!��f��]�ۆ��rgu8��}ߌ���~NJp�P�����^��Ma�]�W`M�?���Ҟ~�Rb�^�z��X���/�w����T����l�{X|:�<�����(�Ry�;M����h7�.9+F����>�]�歱|��'*�v��I�����I}����94�3��i�d.v�2
��q���	T4�XUĚ�`�f�����2NL���t>�Qk�t0�B�c[���+-I��W�aP�#K󸕭\_��z�@��-7��D�Ǚ��ȞXv����B���y�[\�eZM՛��H�Y�;㫁k����X��t5�:���i�%�]Tӫ̈́<��rߴ�{�~�
7��Q�7�r�т�w��_�B�JĐ�8w���u��x˩J�s���j�q����+�BM���C�?��*�G����oʛ:"se���\��@��r	�f=���e�ۻ����v�V`DeH�ExK��2@[���K���d���Y.��ڥt��ԲVʝ&�ј���������ڜ�/OƠ c`]nd�x��fޑ�����y�q���]�o���b'"����B��ގ��ld�$�f�$xS��V�zh1W����(aߵ���Rh�F�Z��ZrGWG���)���#�K0��8
�$�6��wEy)��o�k�(y&x�EU����9���uʻv҃�;���տa؇m��n>�T��a D�i�\��(� ��@iW�u����WD�oƼ?;�+6�N��S�F]�nUW����@s�����O]��'� L2ً���ߦ]�g,�8�o5A���$P�T��Ȑ)z9I�8�l����	���|W�Z
쓧=V�1N�bdF�~��	�����79]Y��T���� $6Ɖ>�LE���g�դ/(W���?Vz�,��P~�=�M~�_�;�9*D n��U��#M���PR:u�≥IO]rV���o�<�z[-�\��&Y/45�,��7�/�(�m�k[{y������Y^�SI�׳��	�]"=�C%�M���s�'ٚ�v R�M�Gu�Vrvƃ���2N,h�E��P|F�\A�t�A��E�}���7j_*P�j��z���9lÛ�Q[Y�Q)�މ�����3�Nj�h*_�/�<�K=�l5l�Z$��z��HL����?�ӂ��S���3^
�*w���7Ģ��z���^����.9,�_�j�C����� ��P;�٨�)���Fׄ�r��Lz���O��2�ݗ�I߹3��fU���r�$陫���z�(��{xXVp�`3*QA@W����3��$IR�HN�$I����4��<���a��}���s]��s�=�������nK����f��'a��pF�{ּ�&f���03rx<�u ��`�oԳ�p���O��z�+)*Δ�>x���Ѵ��W�I �X�g1R}=��9zF=Oi��۷|0�f���|@�iD}�u8� g^0�^OS��`8�HJ�	�������pe�?e�P=��ĺ�����o�h%e�2V��7�$�=꬧�ؙ�>�Y�)��y��H|�*ς�Q����#n�s�hjOE�8�s>[���7�8-_VSX�_�u����65U�16��M�6��f�k݋�j�����"Y�ћ2��_r���Z��5��6�h������,��T~���%�n��(a]U�Tja��f�.�η}f�����T?3æ}�'J�t�� �=<ò*O�Ct�u�Ps:���?8Ѿ��^�ޛv��c�c�	���3e/�>�M/̅����ŉ{�rZ�Z=�Q6sm$vc�5�(`m�2P����1�ٱ� �T{+?�rPm�6}i���)�ĥ_�'\�&�rB��#���o�T9����Ci�����ZފcE�dg�W��sU]qL����a�Ms��@�p* ����k�MWUD�$u���<;7;�ժe�;;�g�vДq�)S������1���E�y�|ѥW�,?��x(�Y���[����|�9��d뛞L�u,�4����tʬ[��ð<N�p�(.��
���I��J�Ȩh��_vM{����3=I��sX��T`P	7��Iˎ�͇<�I�E�����}�S�� X�m���ӉN��]ݿ&����_�5ӡ{4:k�����z�x�5�|8M���:�7v�@�d0��V�ڞ6ۭi%b��G$.�-�Y�Э	�v.9����u�vO���*I�\���,mǪ�1�����(��2���&��G���j�~�	�F��|J�M�9�����l��A	��9�'�����w��,RY4��n�{߶-<���G��z���1���nc$r�Tt�	�9��F�V�5㢰5���_����4m���'H�qŠX�^�.�1�z���gK�I�ǡf 8���׮#����<��ư���P���uQ�Ӳ���'sOm�æ��18�e;	����1(����;k쭛1P�m�دmoi�6�E������8�8�(@��6�V*.q��T#�J����Ǹ�6�_����(7�W����))��q/�%��l��B�������|�s�#�ؚj��蟸ab�$�"�)�������t�*�ܣ���6[[^����o*'%o�k/oׯx������#ʞ�$0ks�Ӡ�IB��66�i̥5���?k��T�����sG�vO����N�����(z}A�R��v{C��O�뱾NУ��^V� ����ņ�t�C�(1�(�4WY�<��cW*
�����6�rQ��qZiz��c;�4��
�מ��� ���ԃ�J�ě�K�@�l|��G0
_�,E�������W��0��
���pm�����`܏C�%�u�镠X����Rps�����t��hVn}l�@��Dg��Ci2[�ffP�~���fl�W��ofҴ�]wRP�r=���|��M�b`���2:��X����_�jr5<���閼���;ZcƊN,|�*L��@~�X�0u2>-��$���ϮF%�i�+�T fm��P�Y�=c��]E�ȷuN0��1|I���f��g�����8�"���μ��</)��ួ�>�[�*�A�Ot<����8���MnFj*D���P3�Bo�������s�X��� r�0��}5�ߢ�xՈW�w��#��j����^�(�]a 6��������e�L��]�FB���E�|��oŜ��	����A�Lo���~��o#3|�QN�i���t�)�+�)�3o��xM\�9��[H�ǉ雂h�E�H��+�=��f�8r�N7$�D�E�(�U��S#�Ds��S�Ⱥ�Քva:��d�S^3���we�V��jC�y�T�n�KWPES�H[*Hې�����68Խ*m�un,�\�SZ� �J��}��pIn�P$⪂rN����C�'Q�Ɏj"�s��Ď,���J�<�b�Z?Vn��5qnU�L�Ꮮ}B�l�]Ĵ������q^pĞ�z>Ɂ�3+2N=�D`.\`$���H��Pp6�9�����Rمe�Q�� �v������?L07��J?�o�Z�������:]�-le�~�Ĕ������yw�R��O�X�{V̯��zy�P�!h�Ʌ�K�� o 7�eڳ�Q��Ƭ��>J�O�4�A�����)��S��9X�f�/ F�H�m�
B��c�l�k�[j�j,�?����oZ�}`����,�H�H�T�u�.J=�J����z���8ORc/s-IN�uUKPCG��ȣ,K����l���4sg�,�TÔH6|���a�|�$��?&A�����O0���t���ӯ�d�K�ڠ��B�*%�8Rp8��IW��+���'��c�e��>�����83eB�G��t�'jϫ�C�L�fZA��;�
�f 
m��}�4|��Q�Lz���;Ysց��Nf�y�sTU�b�w�����㒢B�����#���ܭ��;]f~��6a�:�'���F��TT+%�ޭ.�?EGH�{�K"&>��ªs�k�cRk{�ua��i}/ gk?(Q�e�՗��
x"�_(=̟��~3�41;A���@4&��sz!�+��Y�4Ղ9 ]�5�J��<�R0h5��vJݚ�_ϥO��B�b5<�i��sC�ߛ�r���b�=�a��&_�)8�����+���^ �;�Sb�7~(�_ �\
>Q���i� D��Ȓ<�i���X��r`��&P��TR��.�kɛF�^�2'�w�I��	���~�� ��5 KyM>���V=^�j��!��o�.��#��>"w�f����S'ݝ��J��q�ف�^�/�F�n*k����#|��ə�^{���+���~���!�O�˴������fÌ���iBX�vW�
k�W���;d͸���dV�����:ɕ2*;T,�͟Ng��t��G�B.�w	_�:�13-Z�4~�J۷�1��`&w�����(�A\jXsH��!{�(���}�j�A=���0����O{=�~(�{ZN9��{qn��B;�Ij�
K����	Lp� �o!��D��>��� ��N!M���C��ߨ�+�Q��]�p<��yB"�>��ϊ�(����5��Q�aNET�
p�Ǩ�(��>F�ܼ=7��3V&)���.$c�����R�.<CB��@e�Fkܼ���-`k C��1�T�e�q�M ��Ǿ��`��@���bTqތK���&b�>�:���nz�0�
���cx�����̌�(%M0�M*���\��7�~YWB�F[(Gu�K>v|>�S��T�񣅫�	�e�> uG5{�3zޤ�����䤅�H���b���+���g'��7���^>�'��Kb�k�OP��p�1bpb�l�h�ut�A� ���W���&l��=u-�ٙT.+����3���H�6��A�?����7j��a��O��)wH�����v���wH_�s�e�OP�!�=!1�|�T�+��R횒�y.o0�u�#<��9:
H�7�jހ+Z���e/���ũ]bd�����y��t�3�ވqR�y�5�/�)��gD���o �o��o;hy �K�=� /\��4*��<ؚ��=L�Y��=(7� O;@�\[;���@�����Y罭�r$����J�`@�0̺�K� ��9���>(�U?�!1kd8�[AJ�7WL*%X�X��hFp�~~08��}�oY��]y�u,�w�,�P�%��>��ޱW �ǸҬNI�ŠQZY@Smem6�aͦ��>��AӾB�N�8<	��ʂ�V��3��)6��׶�?#R�u�h5-h}O h�_���<^��/�����Nѓ �����=9����_*����i�Ǡ[�����k���^�q�B�z��IH�N�һ.����<��b.{0��Ye����%6;����i��6��'0m{P��L~��V��-'���߂�������I�J--|��9!qb�|`�� 7��6ٵIܽ��Ӥ_3�PB�E��cr};���B��{�w$}�M���rY�o�a#3�UE[)���䀗�t�΄R�ϱ�8'o'iě;��*v�_����+MwR��E��_(��+g�����-X�0� yr���\����{.��x*wt�����}�Ɠ��p~((�xi���ko���[�����S��4)��!�R���|������A���v���c��d�WXb#	P1�� �ԯ��vE���{fv����|K��DQgOh����y�_؁�y�R�E�VK�(�ԧ�J�1���9�w<��CEw�����D
܀V�߹���G�	��7�R�T�W��1����`"%;��2������8f����)�Wl�,V�,Z�ՇOS\���\����;1�
�����z�H֒�al� 򭐲_���H$%�ڮ�T�\���;����bK��`�� B暈��}��`�i�'e֩9#�f�с'���P�q�is�w�y{T�q��TDy�U�|MmajJ��Ѷg?�l�,��}{�w����B�}�:�j�Ԍ��!ץ6T*tʷ�Q������͝�Z�xM�.ׅ�y�~��zsHAU?�o����.g\�Z�V!�֨�p��i� v�'ײ��)���SoCu���9:��Lm=~A�uw�u�d��{��-Z�~���A�y8��¨�O��6Ew��z|у��Xll���g��F~P�oz�۲����b-�x1B��
(eޥ�;oM$�uvv��N_�/��u�	�����.uG�@n=k�ށ�����#��Ϸ���|8Y���Lv@����bgx�ǈ��.�G�.J��gEG�,��#eLz֣��k��!�K�vne��M���z�=�+�G�
hϯ�w��*�Y��9�
q���M����CM����g�W�w����2Þ���)�
Z�@�>nWo=�&����W����	, �'6�γ�f����W�9u�k?��v*�����������/k:��G��K4�JRv	k��W�oAd޾�i1惰�T��:�W��pݔ���F�����;�k<�C=�����-�N��w�Ue����c^sj&+���'i�xQ[j�l� GWZ�A�!�t�`y��K�5�-\�o O���`���@����5��t S3��/�G�In�-��.4>����[tJc������`ס
>]����/����� ߩ���o���k��ϩD�����K�OQ���K��9h8G�|!
�ݹE!���A�ݼ�/�p_㫸��|���*��-ᕺ�/�?���l���<���7@4ε���ޮ������$8	�矙��?O�����y���$��.��9����mJ�jRF�X�<K��ug��V)�[�9@��mFBM�f1���T�Yҝ�s]�^�m�:��6��6�W�#�|��&?�m��d��T��N���fU��rIu�\'dW뾆�WGvZ�g[S+� �)�I�O7^W�};��\���ڭ"K�Y����=�9�I:`��mEv�3��VͻI=I{���6�+��=J�덫�EԎ�,{��'���� m�����?���0�2��{�sA�&��{��oB�P�(ݙ�"��Vŏ=�/�D�U��������� � �b�����cf��d�fc#'��i��F[Bq/�8�-��3��w�QØ�&CǱqF��c�fOO�K}�Ț��V��<����i/o����:���#�>��+���1�xHf� fWܦ^���B�(h�;I[= ��Ag:�*�v�`^j�٪I!f�o���C-s	���[k��|j�,nP8���u}���ǋ)݂Aݗ�m�|����rv�6�G]�(�*Stv�nl_R,/%o@#L�i����A~l6w��V�����}�w�Lx]�&�;�s�A#�MWz"節?W4|��<v}q�կ=��sР���<AY�Jx1g���	h��12��pP�n�u�>$��4��pjG0���K��{�,�w�����R`f�W��A����mom�"D�'0�h>B��A�H/����^�ꀗ���
��**^�5�⼘���DwC���_�ˈ�!��7h�<�(���їV��ѽ���8\�f��JK�޷����g!���y$�-0�O��w�zǇ}@�
b׌/%Ń��8G��x`�W)Il��ՄLG�/�[`��pŁk2t]0�U�*��v�!	�U�U�@8'M=^�(�}~t�]7��_w���`a��b�@�Wz�͞áu{ �Z���h.�� �?��]���oq}f�K&��I]�m�/[ �S;ሧ+WmU�.|���������7g�b͵zR/�MVs ~3:S2���{u�u�$�o�q�t~p� �ӷ"��D�˙/�I-mqʹr���%�Kr`VՔƕ��=��j�xϋ�!;K�;,��������z���F� g�|���T��>	7�ؚA�A�������|�o�'9P���͑��������h^{��D�<mna	R�8�I�I��v��.|4[Y�ѿ�W����Rq
�Ĉ�����{���=�V/��]Y&WAuK�O����k�H���5<�v��{^���@"Ѻ�i�)�(�<���WKC_W�!߻�|��Ǆ�!?�+�hp(��N��1L��b���'/w6F��.��z�nN>�c�DߐR�sn%�`f;��8s�w�c�A\e>�wE�T���J��jSa���͘�:
c�#i�=���݅ �JV�S�l�糘���ͅ7$�_(����Xj�Z�i����@�+
���%f��	�]LJ�X��B��8s��wH�ǝ�;E
�e����թ	f��Y��"��mN��*�,1�[�ت�5`u;�!���R���oqIe+F��ry�Y˞� Hq���������֤�݃hAu�����ހu�&]�Ke�*t�9vs����ā�ͦ���1\SD67�K��;��ѕJ0�53,�5��Z6���7MV2|��&��k�q.�7�f�DAٯ5 ������E�w�[qQ��^$�k�Pׄ�l��W�.m/
�����[M�z`a�������f��Øk��wLf��1��粐&��T���ou��_��7����z�� |�""�O� 
ڰS����v63�[�!�L���-���VQ�%p}H�_��B��i�ƘA?�:����&�?�;+E%e!c0�@2J��NÝ���Wa ��������|�L.���q�%����ދ!����s������ĖnZ���F妘[�͆���tg��V�z��Ns���0���n��n��[F5��?�k{��w`�c0VyP��.ֺ���fpՊ?%}`�Br0�L1|����ݟ���[�^�Nuk���.�Ʀ0@��
zh���m}'9r��c����@��!����ͼ�>MN�X.�������e�8�n8ǭ>Z����%�f��a)�Su��H���S�:-pr�*A�'&�6�r,ÞՖ36��@��%�:K��������I$�;��ZX狂��ފ���a�!�,���k��EH7���������k�W+b���BMf��Ϭ�Xdp��~t��f�`�X�]����4=M��ᗹ�ޏ<<Tv�����z�{�x�{x3 ڗ�8�P��O�~���z����E�\nn	%�YR"��5��"�.���e��F�ma�+�����������k[e��+�2��J�ꦘ���B��4D�(��m�xЇȄ�>c�V�)���ˤJ/Y��`_�e~���t����6��ÃC��.�8�($⩙��Ӟ-�E��;m{�MW�: Mx����a�A�����a��6=��RB�'��z�ft11�_�]Eb���
����Z3!��B�B�K�ކ$(n\"5���:��x�G.Ɵ�`9+�Yi���&fh�*U"�����VF��z� M:j'���%�`���3�B��i���w䶶&P
I�J���[w�Qt���T ��^%K�T?�)��_�%�Zu��Z��X��6�h���k�&�{��Ȥ���ėX�mO��Z s�Lx���Q��ݞ|I���|�����H:���\ϟ����PhO���v�C�\6l��ᶼ�����˶�����1-��: 8�!���th�{�p�������<;�0�:E@���gǩO�-(��("%�S�q�����425~�9Qr��O� `� �֓�k�գ�y��+������g/s�{�!�ۭ\K���G�i��C���U�X�5&���������Te��|6CC�ݵuO�}�׿�|#�we+@���	�e?� ��5ݖqD�%;Xڛow���2!G�(b��)����<d��t��퓐��`�8���Q���0X~Y�� ,�Z���%��T`�e�:�������B�#�z�����>���:
�H�y���+w�)�So��E)����
sTL��͒X���}K�T7�9����_Ր��V�����X��%�8i��/�E��ں=�!q2K���b=D�۴.��a�A"CI���h3���E`�s��%��ۄ�ض�m��>)�LO�H}E?g��1x�@�	G�X�� ?�iҡ�����g���_ ��v�0���&4�Q _�+�/=�2���aR���Ue�`.Bj0��_��`W1 �5��<Q�F���O��ټ�US�/�C�n� �w@�8���ڳX#���h���PT�PRԂ�E��z#���v�gu��;�`�x��L"3 ��,xw؀:MJ��-������G送�'�욹=������u/�9]�P� 
�6�}Fz�����4Bf+���a��Ǚ�~��㞟4��4b���(+@������K0̕x�c ��ծ9���Z��1is�[ܪFi$�I=y�hEv���^��1�+�B�K6�1�v�{��>��K������C4HIӱ�ZkBjd��B�	��<.J*z�֮ϗ��@!t��^�wB� !���Ӥ�����&����p���c.�3�g ��&G�JcNb� ���񌍺ѨT^ҧ�;%J%�-y����3���v�i68�öo܃IY+��8�W9	��Ic:�K�B+�R�{����þ���Cxz��a��I�m�#�#�U��0x��n��(J��QO�u'*��!PK�a,����rm�?7�|t*-'��!h���[RZ���M�%䚸�&������p���8mW��g��e���Ez@n.<�(��2�f�]�G��t�����퍐��9�"�?�?����`
==�A�T������6��3�tq���^a2 w^�`K��h�����[�����ִo�",Y���wj0�ʤ�1�S7k�@N�PB2����w��7��!.�
K���;셉H꣼�"H��K�;�st�Ğ]��K�g�GǾ�E�D����	�� 8P"W��ٙ����	�Ϫ��_���B�a^�nl1j��-beY��t���H�	D�|`�5�.h�b��@�����}�j�x����<��"-=���(�nL!��>�V�m����i�5�tN46*~�2��.;�x�l\�l`�k�+6�X�Du��"(Xbc91gJL�?MR�V{�
pK��O��ޢ|>�ó�5��'p�C����
�xt|�����J`�T
b&��(�?U�B���f@��;�h�#���$!٫�Tٹ��3���b� \}���ʞ�ZB���'opn!��SPt]�SڬH2Y`2?i��g����/��,_�M�ֽ�������*�������$�Z��!�LQ%��'���>/��D�T��|�����q��KݤoDߋSgv�xO��u�n-<�K/4�ѱ����䃟�����s{s��!e����`a��3�W�^{3to5g 
�W�4��g���-m��"}�Z�/�x�/�S>��UC�3*0��aV��5\ɞxS�IzZX����@�1a�z}���qU�Ge��"��U]��z�n��c�B4f��n�֥��,�DNt���]U��P��]u��y�P�t�L�aq�}���a�7�|���'4�g�j�\�d[I�uY����w�!Q-�z����6L��� �+�~B�����7�Vh�M�|��&�|TJ+�٣�e��O��6���Gy��h��[JZ銂t|��j��]&�#��*MSOᤢ:��F�͏?�V7�:Y�(Ѵp ���k�g����^�������\m��×8�l��������n׵M�
�|mM���n}�����ᚧ ꘴a?)��ў+�K�5Z�K�UA���u��W;]�i��e�2�L��m�Lrp�N�ܮ5�;F��D�
r_��6���m��L���ӛt�߅�_��1���K�a�-��`�	 �q��/35zk�%�S�IଧR+^l4 ��N�9 "|�/=��� �ܬY+�/�Y+u���'��D:�o �um=:��@|}��#ff�¡8�����Dq��d�{6{��
��U���gO�"��O���Q��/�N->�^�\��͆N٢�Y�i [��%�#�={'z���V-��K� 4>پ�)���g�PѥV���ͷ���;��i��Tu��O�QO�L�]��.$�;$=��i��xӶ�u^]:�U{7P�%���8�&���L�MM����f�e�$���܎�-Ӗ����І�^�;�2X_���_ȝ�����r�h����R��x�B0�4����:�ہ���7����J����ȱ��K�0/�]�{Ig�	~#��U[���O;j����!d�I�>,ޘX��$��ל�~��B&������U����w�.�;P�ﻺu�̒_9�`q^�!q��+�W�sxB�R��h�-�F��o�6)���Y~D�� �[-Q|%�z�Ԕ7uf��0��W��U���Gw���va^�'��byeC�����s��@����V�� �=Ȩ�C����_�Ƕ>xL7��2 ��o��k#w�|�(�t�5qD�旉�0�/LSf	e���;�l��jHC���v�5T�y��@�Z����X�V�=^��~?�����x�C���g�v�F>�d�����;r���œ�T_:]v��7ӑi�7'�&��*����K��*��D3��_S@��З��͸� wiGO�yϿ���1���/J<�b��/�Y'���<�t��K-t���Ao��?��&5�Sl��qhV�,k9����������+�F�Q/�� �+;P��!X��:�k��?�_��������N�K�+R���v�
[]4k5�]��G��_C������M
�$��Z����^%Y�1�\h$�D&v�"��u�8U�����_�o8�N��,�0--��F��ϋ���*'�ޏ�Y�Y���u ��Qgf���2.��N+������fP7��yYՎ�D1�#4T񱗠��뽯�%��:4A���[�;IE��L�olQ06ya�����*_1��h�q�[oWW�O5�U�X�7��X�_�M�W��Ҁ�*�BQo2Z��ī|�TS(o2<���t�~p ��\��V�l�X&��xPk{8�E9"�؈E�#3����;Q>�k����,֙�,f�W٣� ����i�3�������Lø\���R����w�ĭ�U��[������m�ѧ"OSJ��h21M��kUop�����'C-�=#��޲�����0sv�K��+�Ĭ��A��l�6ЛԜ��B(aJ�9էg�O*J��(�N<� �Ur B?O ȁ�����-]�9`�-�%���m�lwR��^Q��e0�]�SQ�P@Wg����Z����������x�8���a�_Ո=����o��>�_ā\�^rx�J~ruQ��ƕ�ja��9F`��b��崪�C�9����_
GIT�F�ʱL�E(^e%S�$꩝ͭ�@]���Z=�Ew�c�BBɓ��,��G��i̐���T��Fl��'=?G���ۙ�5{<C�n�oM| �S7Y�x����<�;z�C�Ŭ��$5-�4��*&���P܇|r�!�ԗ� �׈����]�^f���澇�p\T���=ضK^TR�Yk�XW	��̷Y6�j�S4hr�O B>�h K3?z���7\����7��/&�By����i�b@�K���=��WXA�|k=�'՗DzeFF���L��Yy��~R�|��_ -!{9�]��K���_�8*2��]�y��_���h	����9l� ��o�Ț��ݗ������L���~+);7Ru����4}���6tZ��sԙ���|��S;�K(�9o�'���4[7A�J�����S�O��+���j24���^V�hY��|�I���*��x�:���C���m]�֍9h������t��-T�}�3�ʃ���� ��:�m���G��m_�6�o���y�����Z�2��}9�i�I��x�)�1��'���/G7���Xl0��ǯ7��_��L'W�?d��ܒ�)3L���������ӭ�DT�#�|��Cs�4�[,q�4��ȳ#@k\n2愊��, ���D�h.�rK�:�B�T�^��㐿���ً��]@6�s�#d�zǨ�l2H�Ro�Cq�)����n�D0�Z�P�f�����U�����c@�X�9��@�*���'u���R
�3��-����M��:[R���4�!fN�+��M����_��H?���rݒ�U�ɢw^�`�A`HB,g���� �*Iᢔ-o�(w�/Z	�1�'�x�:�3��v��!��5o mI����i����4�^�/W7eE�4A:x��{_���+�n)��f�3��.uViR�r,�ꁤ�Y)������V���#f`��݋<Ĭ�Fr(;:h+ ejTB¤��u�d"�p�c:�w;���Ar��hF�� ���RY�<�V��l������tx� A�Q��#�T�y�/J�;zI7e�j�V�kC�/�OE� �oq��Aq���^N�,J��Q�,'y���4z ��"�;���ֱԉ/� ����o��%ɒ���0�}>���(����{�#z��h�h��]x���!U�{�]�	�T:S������Y�̻f�Z3X�;D�<(e}�r�����_��s��E� ��,��̃^����Ǘ	���xOB��-��!�9�B���ԑ�ר����iW� 4�Xªߪ��h~,i`h�;3M>8m�2d[Q�l��BO��w�&�.�N�N�Dm)ˤR��b��>o�=�[�����b@(:!��M]$�;xx�mv���z�Mw0�������:��I˶����}���JI�
��1��{��Q8����r?���J��HU�j����A:_�'���4w��ُX�uLBIB�T�\�Ş��ϡNz������#&�
�Hԡ�̲�)�s�v[+[++QZC �����B��"�:��[�N� ��ˑrR�cyk%�D����̝����"���X�׆�ɑ2S����8��������'0U~6l�[zgȄ��X���(�����(*[�i��*��M�1�>.2�g{[�~iі�� �53`��nU�^���6F��VJ�q:�7apOKUx��,e6d���PXL*��b�z+OX�%(�x:��"��[�	����M)����/�� �V�g�8�����q�p/�c �o8�J%h�j �����o9��j��e7�Z��w��l��4��-�ݧ���;9��a;(�@)�����yMCxC����'.H�Ev��Q�J�±鄸�R����@�CjLpő��c��[�~�(K���)�4�K�1E	K{wr}-��J���S��!���E���䱍^����������3��H0���VJ���_`c�a)d�T�R��콽��x�����&e���`"/�c��:|��, 8���b��w�;$A�������*Dд�g�ኀ�G),���0�t4Z,b�*��.I[� ���mFg(��j!c55�6}� 0w�exp���cp{��;�Ձ�S-y��������|��O�|��[v��ݗ�����ٽ�\����Խp�p��Ra�m�4��x�����uc�sX���o�Iģ[=S��n-��ʊ�h�8����.�|���0��[{$�`9|_���=���ׇ��,�b�a�
��'N��\��ֻ\��VX�U;����pi�5L̴���j�3����=5� s	��e/'Ε�%X��y��m� ��l�l鬨Hu�U�{W6���8�l��۟�w����q�D��mۡ�g�_{��}��l�c�c��`������*=ʝP���ъe����Oڰמ�z��V�r�?ͯEk�>j%���ܨo6?ܚ(O�"���b�!�_;�qP�=�K��.�{lMIS����B������`�hy���j�a
85�T���v�Ϊ�rt���簐����BCk�2wG�����e���{	�-�a�1�����e����G�?���;&� k��š���]�jڍ�3L%-.W�(<ǒ�|r��ܨW����;��d@�rѫ~�M���W3B��-�կo��=��	C��F��J�kk	tȚYW|�G!%�������]�ɟ�C�\9aʠ�l�s����JTm��G�[���"
d�[:?��C��B[XyOșjDJ�M��ؖU�2�*�!����ϙ�m�|�d"1����!Q�!k2�$$Y�owL'[ ����ŧ`XP������Q�?�d���_�g@B���=�X�lF��f׵w�q�W�(=G�� !�d�J2��
}��s��!��������rM�`[�_���r�έ�L��"���n�n� ,�z�X�%�$�F�58��N1+ ���o�Evq��Ӱ�X�@�U�w5��UǍ�z*�W�C'5�[�D����}S������]�=���XWN�I��2�>'fv�̇����W�כH��A�ߕw�9��⏞�Y�����/v�%��EnT������!���(�BP��S���HҍAZ-�����d�����J��u �w=���P�[���Xu��5e��&,/�[�O>�,�SO�! ��4�]�p`x��rp#F�}�y���L��4r�Ktj����)��U�I�y��$�d��w��E�+����e���~>@��x ������a��uǱԔ��~�l��w�0����F אI�����$&+�vN����w#p���{�v;���۹����}V�L�;~��-$]���BǮ�5%|v���Ξ���]_=��?dֿD�����0tʹ/.l�/&+���}[�q�`.�J0L�G�4_��k�l��k>����;���o�$���
:�$�ǧ���k'!sa�Q�V�>$zp���d����DeomA�8�'������F���N3����̐3R�c���7|���Ɯ��wv��#���9s���A����`��Gމ���&�+`)�27ko݉h���%=�Qp][}�<�z˼���濡D�y�qy�3 W��~w7��~q0m�Z�&��L宆vqtF_<q�M)�˴ܾ{VypOx�ҭe_*���Y�Pk*d�Ȼ�C�{�����"�4ծ�b��6��s� �gΏLf�Ē��������Y?��`��馿[������1>����C�%�C�x�ӽ.�a�t*"���t�����y�A���d��Q4r���l�)X'F^q�)�\�Ǭs�LTT���ԩ�Em�ڐ���z1�o	��f;Lqm�E�.���<1`֥76= �!8��s =�bY�ڴ����g�D�,;""�6��4�����C��z�F���k�9���\�`ܛY*y�,aw�[�K%��y���u���q|�m~L$Av��*�ܧ}G�ύ"�X�>!�����W4[��xL��ub�B-����%6᮷@�����Q��G��OO���!�ę�X�l�S��.(z�9�����q��Lp�%�V=J������B��-M2y�|�k�(�1�O�e�m�2��$���A�҉X�+���b}@�f>� EKz#7�v��| rh��M��"��0�g�'{���X����l�庫t���P�㟾�4Y�����|����@��w�)�ח��vݱĠ{��4�4�lNS.���Ԧ�a�;NCs/|9���������1�Y��|z��`/��2}�����	�m��H�$�!|{���	 �lÂ˺Yt�"�&��M��qP?�gr2C&jիA)L����2$�rn�A���j�3F�G��9U�� ?Wx��P)�F�+'�p5�����?�m��h�$�K����XS��shqXe�[5�6vcҬ�r����ږM��k��~�*�@���YYq�닾 �Q��G0�&�'9��m��J���)�k�l�m��g{;���@".��5N6-�}�Oi�@v�iE�-��!�<O�4������1ˡ�-*��c���|��c,��^��!�X{S��ior�6����e��l"5��w�� �b5���p�L�f��`�O^Y_x�g�jЙ������ۋ���"��wfn����HFV}��AapeJ�a:΁��6������A�ܴ���c':�a�#��������PakȤS)j4�Ю������҆3|� K�fju��T�\��2��N�����������f�����"�OW�G�W����a���zѨ��Q�4�^�3�	��a�n��A�mm�iD�u E�!��z�|ri�r`v
�?{Xy;^����/��b�eb�O��ȹ'�w�ז��$���_9}�U�#|:>���!��� w��|n�2\�E����1��7�n��#m@"<@"ȉ8�'�/'����U ��+��������;�P��#�R�}��-(��+�����*�H����I���ݞ
5 
n�e�붯}IL&XV,3�y2�㼫�4�Z��#���#_�f>��;6�z�.�,�^+m��z��7ٌ&���0��yk�=���(�����؁gC��d���U�_�E�O @q�DӲ]��X_�� ؠ-2����#��4Ķ�"?���\bl��/��"���s����Mg�'�|��{�����:� �7l?_%�O�!}d�n�!�!!�	��4߾�,�6�E�M\g	�D5�I�1�������-�e71*%�������8R�� ?%�3T��|�Y{f�bhG"��Iۤu&������o���s����1�Yl�4^."E��WQ 	]�@UI(��Zq��K��t(�]�?��[ ������8r�+��g/�9%"Z'�϶O�~��:dZ�!�Ds=��靆��\����y��<��(�(�����fd}�b�����d�sQ/�2�j֔w���=���kn�1yt�p��)��N�\u�ABU�c�0]�CVi��U	�����ݩE����B���!MS�^ [�$�u(]_n8�����x��+��1Y�?�m�ҕ����k�z�p�5�L�c���w�����uJS1T�����D ��q��L{������ТQt]��Q�2�ɗ����4��F����料3�:�%��Rg�n%}�(�#	�u#ߍ�������j��O`�.�'� �	��RX�4��-��d��I�##�[���VSv��n�J������`�ik ��hL)kJ^�����d��=i�84��b�O��ǀv��б�P~bG����dǙ��Sg��fD��mZ�jXz��h�S�7�T��� ��ͼ�QY��WL<���V�&�²�a��t	.�e9�DѺ4�:07�j��w�q�o��l
ߐ��=����7���g��K���nW@R4ͨ��7R�ͻ�����:s�^-.K'n %�!�]3�ɣ�ߊ�q�4�3���|�~?�����R%��o�����R�����?.�(}�ڢ����m�4w����zۏH��B������5~�c�߻y d�cK6Ba_L�7^�n-l�����`{��}���1G����-r�~���Oܚ���S

��cF�X�H�E]�v�3و���#ː#y�A����@�s�ډ�JpJ��B��L5t�q��w�MK$*&��Ҋ�`�rփ��V�d����*z
���> M��&��߼�A=y�I�>�ewuL�I�Q�16��D8����Cd��r���b4�J�5�h�Ͽ�_��e��a���x� �Z�J��,�D��0��A����&z��=�պ=�kށ���:�Z�C��~!{��Ao�}���kz�q6�ٳ��88Y)I$t�I�?=7�X� �U�tz��p�
5�1�=�x|��k�k ��㓽s�L��{��E��뮸�]�iE�`@@� .""�  ŀ Y`$�₂��U�̐$QP� HΒs򯪻q��u=o��?�:5]U���>�9�ӥi�Gk�"�?�[��ց����)�]�����a�;� r�����i���"�����޴�Xl���`��m�@}�(x�%6�2�����c�����F�¤M���M?�M�Bp�	���r���� ������V���;G��-�5��l�u�J+kPڵ'X�uGFIjߎp�XZ�T�TAlf�[����1�j�&'*s #����܊d9���m82e����b�س��*� r�8�1�),��FӾ6�e,��w���1;?�-a�:{,���e�C_�[���C�/��Ye�����i�O�;�og����p�t��(,gV7�!ԭJ��s6���.�0������y�M�h�!�}��|MOt�LGbï��c���j~��1�ĳX�����z�}��Т���x�aB5��
F�;�~���S�����/�R�BL�+Ua��^W�NlѼ"B&��Z {*/�\��M�M·;�9� �v�V��q$R �K-J�o1�� ��v�۶K	���z�����Ά!�G�+ف��y�_���8�����o�����*X�|&þ��جΥ��}+�h�ZJ~!�xڄ)�-�/��:
���)�!`1{�u9�٧z!zCX[��c��V�R��x�ڰd���U�P����&���ry�᎝�@�A�"��hf���9��.���Y/���`����$�Juگ�/a�d ٻ�w^t�	�|��&vH�S��A�޻AldE��_���q�0|��|߻n@���M�ⵯ�xJ��⁂���r�o�X�)H���F>���8hMt&�ӿ���ۡC�V*��m_�[�d�K�R���6�;/���Z���י�Cl�����FS)�ZB#'�\�ָ�f׏��1� �w<k�=��q�(�"e��|�X>�	����O���D�T���툴�.���D�������2�j#�@��o��!B��z��N�ހ�˥�,A�)@4����s�/�X��*ܹ£K�p�b�R�,����TJV0'�x�Hk�ol�w�qY��
`%�)�";��e��\�ǌaK�
�׼G��/Q{��L)g�.�u��~.��o���#������&�iTZ'=�=�x$��$�v�m�(ǰ� FM��s`|��q2�A��m�M����HM���bam�dk��|��[�%v[ß���Q����o%�컗�,M��c�;(�l�M�MG�d̪O�;�ZQ�G7m-�l���K�c��)�>k�Z�����)w@>�����=�	��{`ѭ�&è�Kzo]�k��|-�e%\g}��}̡Je�^R,�M��,R_�=&�r���ĝ�����/�"��Q�U�6c�4x�©�팿A�����C���A��M����+�x%��6ੲ�hn�F\��y�O��b?g��N�a>ݲ�{E���~|�������CL�&�4(-H�l��_�M[Y86p�����:�Jb�5�a�p�-}m�nL�{0�v9���_�jf���6���-R>9b���>w��O3�O���@#��,��3e#L����l���ZP 8ht��QȈ�I�7@����ҕ�A~�A��J����,���Kej���PJhilk�����Wt]~L�l@�1��e/����b@j�J�L�N��8���S�)�Xk ~�� 
�W����cX�tyG�������dR����)x�œ���V�<��&�E+�M�@������S��Д�m�ࠆ#f����\���C��7U ��2XJX2�1�]�섽�<�X��XJ�������H�ϥ�pཱྀ�O��уR^Kԁ*?�<������ �xi��!�q����������&���/5).�x�O9c��~�]&0]��J�o�#�����{Fd��J��Oc'�@D�j� �F��{<�.ƙ�X���E8QE��T^j����m[��,�ZQ L+�UK��A�X�>˒E�Ya�Z�ne��
aw��%��YI��2�CT���\�Or!s�����ۍ�@�{l+'��\����,zC:��z&q��?R�қ������(/���XTfZ�N|����%�xU	(u��-h?/;��� ��c2�!rM��~����Lx����3�=��������6���ͦP�� ��(�]��jbܙ�݆0̧(�E�&��[�*���y�����aK#'(h'z\�73�0cs��G`0t��Y:��S��~CL$,��RȔ�^����G&��z�Ԕ'nVZ2��niT��U�v��&��*� �#O=!�o����c������׎
� M�e/T�tI�n�N=��:�~�Y'�����}��c'���(O5Y�;��D"kk�����S9[q�
?3Z�H����7j�b��}�e�7��#S�R���K�7����և�g�C��r��
 ���������`W��9��Pҁ���bsk¹��-�lRx�cv��#��L�����OY��æ/����l:Qmz뚓��B�o]j��U�6+zq��|��W�<0<��m��$�3R����	��쐢��?���ڷB��j��9 ?� �!"]Ʌ�Cn��p��%��e�KBAs��cD����nc���� ̐�	;��ݝ�j�H�Ch��@%���J�l� &�H�ܴ����i�gj!r���J�
Z��2s�[�N-B)����|�e�N.�w_	�%�+Ͽ`q�I�Z�e��_`�J���D�^}���ȯ��nkPY�nV��m�d>V��n�n36�����N.�=@M�����ޘFl:�&�BX
p^�>"ŠN����	���L�^�R�Y��<@^��H���oT����6K|�=�xʹ��l	F:�1~���",�G�g+��ȝ�0��=�����k#�U�T'��^��s:Ժ���U�� �N�T#ʚ{9��&RC�������Î�Y ���[#z�Zb6���[�5�����co���w�6<�`���uE�i���`RL��	���}�%�ݺ���� ����ODB�;��[��ͪ�����Kh�h�ws!�t�ZK�_�p��4GՓ�b&�&$�L1�rB]��T��f�{a}R	Y��6�n��1��A��gw�y�A��?!Ƽ~Z?�c�Ύ$�Uկ�����(@E��YAE��,�j>�[���g��KQ�%#�Q��_�a�I|~R4�0#�M�~?�F�.w�.�?�F9yU�A�y�%Vxze�+oY8/�y* ��n��G��;v�܍A����X���L�漜:T(4"�k��o�\���$w�~��2�}��|�M=���| �u��Μ�Y&y��VD�&��W�����O*c=y����{��Q���$��:ӐM,��8��k�m��h/e|���n�K�*b8e����-:L_qAE�5�4,��j��K�7�N�Q���m���H{��P�M���?�v"}��f*�Hl�Mϥ)����P�P��3�7�pB��:�,�#�E^g+6[jϸ�}���]�|v������/؟�<�T�����uK�x:&>�٣��YLP��R���eS�Y�`���A�X��L�jn����4�r�!\B����A�Z�m��,G}�k#�4c�f�i>�E#��W,3O	�Su����I��o��@�i���z.�uO�r�C�QG���0c��9🭒.\�����5�UG���ɨ1Gޗ<u�g4�@K]��<Z,-�eW��/�-���ǫI$��c��J�<�6�O0�nzq��_����T�U��ѓ9�Մ�n�O{�e���}�A�����Zb����ǡ����H�n�p�v7�=�~�ȧ�ϴp�%ԭd�z8x�E<w���_CJ��Õ�W]|͞�}�l��������>!�n�Jw�L3��n�]C�gʍe�W�,$��C8q��x�`=��ĔB~��(lX�2�����}������>�߇�������}������߇w��&Rnh͔n�_��IV�{��Kg��b���O��U�wM�7fM��ow\�tڞN�(1��V�r��Jz<Z�����k��+��k0��a,�A4k]��&G�� Nk�>{t�C�V:�gyA3�#}ETv����f����ؽV�}o���^J�RS=4����[̽�7�3>veJp�S�TM�t�.8[����f�A�2I�q�н�IU�2�+7W��%�ɌoVʳ,��//t^I��6�6?�>#������4���6�ʧ���?�V����L���cr�-�}iO/]�L��ط�����<|=j���S��RB�=V�`�����9wbO)���a����o��������$��G�0�J��O���g�v��y������ �, ��\;$�C\"U���rj�	�,N�?`'�5f3,��.şX������R�7���^�;�Bh[�{�S�ŏ�p����y�^���zU���_��8[��~�m�m���Z.b��cǿjpGr'Iڼ��h���0X.7�Z}��fn����ޝ4�J\|j�"�#*az�+9�\Ò�y��vM�&�ZW�j�l_,p	�Noۦ��oyf;���t�Һ����N�^��0��_bʵ������il�>Z\t�'���h��ө.�tO�z%�H�
p�d.�B�z]K��#Yo�ɩr�h�ҎBKJd
�Q���e�,M��=�[�3,���F��ќ�g����"�x0��위_��^�O+�7oڌY;A�^��F%#wv��.�`�ǹ|�7��v� 1�Gu5͚�Ф�}��2K�J����"u�PO���#�Lv ;�"S0n<a�Ԗ���Xӹ{��P�d]���kp�MaW��,�Ľ�����u��[(��Mر�7D�I>K_�y&/���c�j�q+�OF���Iuqj^��A_��5�lXa�CZ�dh[݂n�	�`�5�$��L=���H��/-22�K����+Nݶx����8_�5�.r��=��nh�_1�6~�N���w�P3��*�?��p�2�8�a�#wMU���m�L��p*�mwﬠ0�0[��yib��a�j���4��8��L��v4�4�^���X��m5=�$t��13�^�~�o07��7�k�}���y��]���l�,Z�u&�o6�&ee����>ʒՊ��V����r.�Cm��_g�{%F�g���32l��u[���'������C���j\���%��X���3lZ/�n^�uIzhV#�\����*Bcm;�4ܸ��Z_|6���,�|�䎷�)��`"נoIQ�b��6ȿU�1�C�ں���~'��BЯ; ƙ���[��9�%�a���ř1�L���_���}i���18v�_�e�\-Y*_<�;���oj��a���r��ݕ^�e�M���I��n��q�:�#l�>,5�W Y8��挡Q�9�>��_����u�Ƹܻ����q���sM�$�2|�.����Q���w�bNR��7�Du�Ǽ��z?Z�l�(ꕵ2���lޔ!<���R�H@l�)WW{��	|m��y��FZA�dn�K��pi�<h
3>��v�������+ղ�}ߡ�T����c�ϑ�֐S(nmVHjN)ƫ����b��m��vJT2+� /��&�k�8��7)S��[�\�a���4�[�����lm]l��6�<�zr�X�x����x�m��Ya��Y���QMN7�V��s�t gmHM�@�xJz4��m��G#4�����HC��FG����ik_=z��������낦[<�uZ;WÉ�&�96��H�TZ�t2�j�m�)�� �����}�#�"�����^?�=�̍�ʍ��[�qi�8o�r�·�P��w9�	k���Ԍ �Ѹ4|]`k�lu��ۋ����%f��YSL�y��;ȑn�q9}=������1��}��� �Uk���q��-���)��<;�����/6�'�����h�gId�۝,�_����Tb}��&�]^uC&�4�����©Ǒ&7�c�����9��V1��חT�tN���c� >�й��&?ߨZ��)���G�nd�,�����'���/z��Rh~��R��M��������o���	�նj�qF�MRՑ���Z��vi2�Wejx�*������ :�{���=E��[�ήܚ��'}�D���Ԙ6;�L33̽��1Wh�څ�ݶ|���\�`^n����!e{h�Z@"�'!B��H�B�C�0����I�cT׌cъx�{l�k�
R�<��sP� pj�w|ݧo��$=�_TTy��c06�.k�%��G�Ͳ����\?�H��,:|���9[59��/�5�w7����)oSeL�פ޸fK�c�6wߟ l�a�j��V����?�a�p�9��Sd���R��׌R� �j3�0�ܙ�/i:�L�� /�l�X�:�h�ɇG��9������t�믿�Z�L��-��c�[U��}�<1�G�<����\-ێ= �-�s��QI�a2d](G����7����N���M�rJ�g��� J�ހ��4#n4d�H)�m�q�����A�D<�s! HB��L_�hӉ&!~z&�TԍE�lq^󣒓��΍74%;R�Ǡ�k6t��gMέ��k?��a�� �R��SMVX�ä�د��f�!��b��B�֑��Iʛ4�xf��)��������[᫦%��[���H�@5��S9x"���x�uk��7�D;ܼ�S�u�����$�&���������j!�.�@q�(�Mp	m1=� �A�m��W��^0�W�m��&�1m<�;�+��/��˄�] �;�������H��4ܑ���y`wN�/J��yyf~�[/(2U�Q���~��[j��ЉOx�l�ι�ݷgj���/�(�I~)tnq��w��y�Rf,���İ`���5���ݘ��uN�"�Ó�u�L��L��r�w;&G]��5}�Ѝ��Hl�0l�O���_,���H�T�r��S�7A���͏W��ރ�V˝�_fb�uhx�!���*,���D�Fɘ̤���X�9Ob�O�fY�y_��?/�h}3�*�r�=�8��J��^�_ev��͘���y�u��?���v�@O�|�p��Ə�\M������:�m�-�W7I�6��`l\T�n�:�4�rWx���P�Xl;*�Ĭ(�����=�����LlK+������� j��ݩ��7�-]}@��h����+gx�2JڍS�P��4��:o�ju�oB��d�aoF�N�n��V���ߦ�>�l�=�^�W���3'�>�40�����K�U<��m�ٱL�s� �wӲ�WI�r�/,��ıT�[TA��5g9!�)v˳i����R��N�6p_ �'N�դ��x����ϔ��M��
se�]�^d�y�	�	��e����m��c�yw�����A#k�7IJ`��/�����k��^U���9)սyST�Y7��.��J�s"�.N���� Z�ĭl��"��&�A�^��ç�9����盜wv���ݚt� P6-M�s9�������r3���_���������m&ҙV�w�.����B��m����٧WV+m���M��!ϭ2\q��@�v�1�Ⴎ
�43s�O=��|Y�[�������+�g{��\Y�����
�v�+� >�8r@V5'�a@*��.��s�ƚz�����dZ��j�Tz���/�4��L�����(6���x	��5���Y��2�=����r������±�'�w�W�� y�ܼϻP&{�Z���l�U����� ~�EB�˩����fh8�+a+(��Q.����VJ���C����_I#��4�}?	����,A��ͅ��,=��ձ�t��2��Ykt�zCɶ�P�:��6�Y�9��`�jz��/f��Y�nFX��J�	��Ǔy�λ@(��$ ��)�����m���"�?PrKٷ�;||��9��-.��^��&B��$����s%�����'��V�ra���� �R�$�q�M�:�,:��;�b9�\K��i1R�������Qg�	a�Rj�ə\�K8[��o���n �X��ej|NCQ^N]Oy�Rx�[����7%���P����+)!�?�0�{GWI���$������e�eZ#��#���9��^��ƴ.q�1'����^�h��m���]����z?n��ޝ��-Ե����>S���)�m{�ȝ1}����	�,b������-Ԗ���c��__�ʘg5���Lf8\a9��6N���k_q�CzI��8�I���""�`pj�\+D_o�����������E̸2?�[���D��fC
��b*��+�<X .�\�5P�:���O�S���oj�T�r=0U��>�+���0�nEi#݆��h�_й��=����;9�)�QS9gr-�|.���u�ѳ�j݋��tu5t�i|��ƮhI%�I*L�s�s��g�9yb)`ƣ�����GA���r�A�`Ͳ���{��Z't����p���/�	_�6֧Yav$1�@�:��-�V�8v�M�1Չ��(P qn�]�?݀^{����1K	*h��`�����$�
���yS{�^��u�T!�5�S��UK��:��[R���ή~ �dL_)j���{�Bi��[q���?�8����R���?ٕ�CKb斃?똈�,iđ����s�)������k�l�a��=��"nN,]�eZ~#��C�!��F��p�1@#�M�r�����I���������BRϮ�j{DBE����e_���e����h�u2�P���Q��
��=��G�d����{5��!ݲ#���YݒR�Қ_�/�b_���?��#��&���
��RSWcb���F�G�����L����.[e�n\�/Y7�Z�?���=w-�u��~��RB���R��G�5�z�HW׬�:�ʥ'1���Iᖫ ��Mɏ���g��=!�Bl���~��OӍ�H�Փ��>�=�q	��ܿޘl�'�C2�֢d?�N�p�Ǔ�����4m�οhu����~�
j0�,F�)����'gt]A�<�B6��\eU�6�1v @�~�����v�:	�ϝ{��!\";��'p�ΥQ:kA�[�{��ʈD��������x`Zݛ�Ni!�-��50�Gx���N�y���_+����%�o[$3���P�����0��h��8�c�����f� ݖ8�74���`{��g�Ǉ��Z����6��g��C��Ԕ�ICkPx)iȬ���y����axK�d�	��{�M}1 ��Ĕ�\M�#s�_?�~ez��s��C,q�j���K�2�prR\�k��̹"|9��NZ@�PO�����!�?��:��?���ӂ5
i�HZ�{���c<j�Fx�WA���1�]�9��D�ˠ��jo+�u�^�������O�v�aZ�����P&�zAZ��l%=	���x =�Q_m�ǔ]%��ߖߦ�c<��Ah)��-7��M�>^�#�?���+E�W+��Y.�R�5����s�T��UyDUI��T�t5n��0)T]��
E����Q
�o�p���/S����� 1:�Y�\_#A��2��[�%�;K��@�p�����r��#TV?��!��������@J�q���?2'�U��:�L�J
N���a}�b�Jcc"B^�Q�/ܐF���+cި����{x<�XL�V��#!�I\�������0s����=����a�٢P����Ǐ`[�CO���,���FY�(�y��ۛk	�1F�ɑO�N����#Jv����+�3��m%s��#R��<�⚋9K����������U��ofq���߉?LK*���K�ϑxQ���D�h��L���ui��]�#-"��d^�e�~�D��۾I��b%�G��.�+8�ߪ�Ƌ�3bq��<܁�\�0imw�!"I�ÄI�0�u��.A����u���C�� ��Q�?8Q����$Bw��:p=K?�iW]@��mq�B��A����F3s}et-G�ú`T�g�l5��j@�tw�M��
�J?�yh��Y�rGF�:�]@pGC��Zo�,��0�,��a@b|�p8RwR��aT�W~o�>>��@�ړ����uS��J~��M8&w��+~��?�p�;�t�h,lT���t Ը*BOR����;�C�AY�����ʘ�X�[�nX��p�@2Zm��W�S�3�ͷM�. �Ø���	�s.��)��CZ)i�9���5�f�D���F"��c����ŋ��~.�Hs��2b�b�!͑�����l8�`=��+����*`^�#��o�.tz�����m�Lm<{-a����J�iKL���%���'�/�g�=jP�"��1��(�Y�lm8�E�罀�ĳ `"��tR�٦�{�b�It�\B�]m��߿[�q?�ǲܲ��z�W.�� ��,�\ind�%"��W(zAC�B���܎m�����¢�;H����V�h�������Ѷ}��'���c���m�&Ps�����Z��Ыj$o��Jb.��N˖a��zp':������ˋٞD��7���3b斜�+1��Æ6�0q�V/Ag�L-]ꔇ��^Hc�}u��mi�v�u?� ɕ0�nȻ0�(
^��*�m4Y��BPY2��bDЎH,B���RJ�5&�X�Nb:!�{_�|@�'�@Q����B
��Lb���Y)=�;Ψ����@��y��b���Ao��f�{��ό��	�k� �k��g����)j�YCƇ�h�'t���ɫ��\P�䤅�Z�精	�'s��$�&TF�Y��R؅����`*=��Z7<	?�ڟX��N�����.����G��%�7"��ǐCV�X��M�ʠ��(o��F����[ �3�#��t�7%�b� ���zAm])�;�;p�"eK�9�E�| �� [������K��>����ɟj:��5�X< ���F��r���b�ϕ)�A��0�q��J�&�#��
?L��Ϯ�㳮gl�|[t��2�������ϦY�ƛ�L�Bn�dV8�0�X�'�	w���V��F��a?u����K��	&�?;���!T�� &�CD	�겆�Oi��0�۲�D�� +W!�ҋ��v�D^��}W9�FRl�!����W��[VLv`lII�2�,^�V=�yJ�k�g2V���L��woF� .��+�ͪ�a���}v>�H�^�����=��?ƛSeB��w���GMZx~| �{�����D/��{�h��v�\�_�2'�{Т��oXu��j0��a� �#k-x����7��Q*�����(o�C,&%���n^H���,˄���>7�=1�;��$�J� )!����O\�G�C�xo�ƱcJ$�<uC�����VB�k�����S;�@�@����In�v9訟�<)�9}�޲r�g)�kG$�şX�;�j\\�6K����d|��я�'�8�4�peO�S��ߢ&q���I��O�G\ѝ���}�l��_p/��H�O��/�Z4��(�x�tn��`�'{<�/7��W�e�t�*4t"�D�����<�01:!��G
R�z>��ȼ�\x�h!�a
��u�K}�d���ƚ.����ܡ�}aK$$��~���L!��L�?��=V��x`���D��:,�+1�+D�Ê����I�<;��caN������(��7�Ԛ*��F���.�R@����D��,J\��2N�^$b��e�s��ɚ��K�ͽ8�;�p>Կ�ၩ��( �f���sm�+2WB���WC��W�4��)J�&�� �ڋu��.�c7�����0R��:�|d�L2������ �wm��}��E
7ܙ�#������������!�O��e,��b����CK��yc�`*b2�!z{�����@�6���/��m0��A����՗�y��Z^��Ⲣ��ϝ�\n�<r�)2q��^��)�a�5�V T�ܜ6�)�C�(��Mb!lw!?U�r	8?k�#��	�=����>��r��kU����Q�Z�g{Բ��[�x�]v=:�bD��ҹU<�����7���c�rɕ`��{ȜY�B�ܰ`N�_pHCs��&a�X���ER�0��i�P��A�sH� :m砵M��$2��W{�1�j�nz�?������������P;��ϪJ$���;����W`��Ӣ���Q���0���RƩ�R�$�\k&�;dr� �%�=l\+����&X�.$�F"P�s�*D)��}1����&�r��˩�9������	�����b�D�b���4�c-5"H���_�M�q�&
��k��7	�����~��Ab ޏ|> �)j�0�����C@r|��D�^'�;P(b� ��?ݾpۂ.��t�zn�:�rd����R��dH��Ȯ8ul����������5�j��>�?m���N�_B�ٽ}���!ma��OE%
M7��j7!�]J�m�t0P�[�%��T� BG_��Z�M�+�I�D���F��&��ԼcZ䛸(�1J"_&F<��,��r�N�O�Kao��-Ý4���?��5|�<B���a��xS�g�����9��/M[���f��U�mڌXn��GY���׈���k����L�/�~k�(���w	r�Dδ�4P�U9���	����i��Uo��T�������#��b�����<��&�`�Fѯ�]����-|��q6��J�Ԍd*&Z���"�r
'����$���ɦ�σ0D���d�GM���"d�_�`�-��%�a�*7%�\n�iɔLW��� g��AL$a����294٫���%;?x�Ʉ^b��X�}��@��d;~WW#/	Ӱ�JV�;�r�3�J����Y�`n�
�$��
�DX�'~,��É��>�ҤK��%�e��A<_���.	X�@�q��
��#����k���`�qph^j1䦠������绸#5�x,a����)����{�[�qj��C�߫�d�����\ż0
���Ejv'���b�Ȍ�*�����x��L=|�[�8xD�=B���׍�c.sq��xG����e�]X˔��_�����2�@�sd��%���Ǽ� .�3O?�/��J�ﭪ�,�ݦ[�~��+5����8�b�U
�E=�$j'c�h@�B`-|+�r�kq�[l��#ۿ<�_������"���ͪ�ck�XӇ�6�G�^at�;���OT���,��KO�������Y�I{x�/B�R@~b�K82�W!gL�/I�ו:%�IO;�Ȯjg���/�70�^(�ͩ
{���z�7Ӽ/߫��m/�_�92�i���cý���m��V���q�k�&Վq��Z!�R�ڗ��[)o_g�����ez�ԛb�]��+��v�s)swv�5��q�d�ZY��P�ԭ��6,�
���z!;"��sl�⑌:������,V.h���s��->�V\�뭹�8͸	�����♅kӵ��)�Z{�##�&sii���p���X�n��X��5�pA��M��0>i��ʬ�d1�e�s,���\V��g��[��U�l-���/�4��FgLS4ѵ�QU���Kvd���EڬI��g(���.ɏ��J\���p��Y�tlؼ�џ���:������\]��CMuVj�[���g8D���bV�#0��o�#���v�Am߿��B��i�����J� ԬLp�%�!�955_� ��״��_���ްG��l�>�w���f?a�S�ݔ��䛌����ڂr����K6_�/�eC�������;\�'�FV4ί`X�.�&�H�	l|Р��}�R !rY��[������P�ȧPk���*�����S�Ғp7=�9�{���ˍ�yOf�zFSs�{�i�LFG�\眇���S�	[gQ���¤\w"����3�Tǎ�[�	/���H�G��|j��P�|��?KI'�z)f�5�(~4�����{f~[D+;�Q?���)���YD����&3e����y�C��%eU�9�q=2Y��O�iM�f�y�5���̠���nB��/0́�܋q�pR���t+7R�EAgO-v���}m�Bg�|7 �"���GRhe���C��lv]�90B#Pf�@��v�+3��`�ߐ��B���������!�C�\7Oa��Xz�{���O�+UУ9x�|N���	��V����l�os{�WŎ�}�
U�;R�lN�Tu6�ǛBw���$8�X�	�SL(�a��="}	ڽy�Be�E`G����4�ФɨT˥����-cm~���X~~qR�ͻmOqu�R�S�/�Ew2Tʉ����8{�Lt��i�w{X\֍�(�:Ư�/i�Մ�/�MlF�E.�5�F�0�h�/����;����*����MvRc�c�N�OU�� ����n���)�Z_j�q�2�jͪ��TKd]�e����tJs�i�_I9/:"a=]�M0�G`��{�'����^����O�>V���
��(c,1]-'b��s�W,�d���_���a2�q�>�^s������
7X+����&�5�:��eW�B��_�J{�˶9���4.8��-�g
G3��d�y��;�Uz�:~�n�]},�G?�<���H�f�����,M_s��U���>u[B&�������=���i;��k��6]u���)�ջ�l�X5�ݹ�pu誱�b�;l�y��gD��<t���?x<����꺧1���>A� �5�4#�V�ط,��.��xE��XFM[ް޽Ŧ��y��C�����k�u�eLs�һ��r
���x'���^��fq~p�f���Ma�X�:��:���KhNmb������=�}tsݡn�
����ߏK�7}���ԇ��?���A~��|e�����C7X�ikWl��������hW�������{�Aj�m��zx^7tnR,~��a����Z��N38j6)�;�56p�S�,+7��b�ji���wy8��9~9��n�w[��D��id����O�)�n��jޗh����4i\XO� �������&�
�Y�����x�Y��8Aw�u���a��NPW�L1�n���8�Vڧ����>�D
��3/�^0�
9q�x�\���]����9���`�)�29K\զ#q�>.ne٨Ñ�7���I�Vs!j��z�v]~����A�p�XU~��� b|�Aih�g�ӌ��{m64�s�5/���,�����]��b�{;�6��{5=q^rQ��K_�-�3#�^�/�Z��PM!�/U?�u��"Ͻ�'�n�2��r<�e�R?Ԝ9b'k
��ճ�м�m�Ӣ�G�[�H[��bw0z��n���)v�M֫EۧT�&�7\�ʞ:T0�v���rs��u�%��|�2=4��y���3[i���t��;ÉO�k^�N�9N��S��R�|��5&������͋4	��d�R!Sv���������g���mz�o�gʐ�MbӴdSD�?�_����A�:��ڝS��3�����8�<�A��Ow���D��*�����p����;�Yy��<U{�~�c�d�!��9��cҽ�d�)=F��!-c�{;/�ջ:���49��� T�[o���eSÅ�zǙ�a� �U�ѱF\��I �4ިZ(}�"Llz/�Ȓ"[��н��S�TvM�g���wS�:��B*�w�.=�d���$JK�~+!��� 0�+�m����7�/h�G��u�������e������N)΢��A5(�E��Ŋ�L^��h<��I;�x`םG��;��f�|R�	�pbo8ߝ}���l��m�URvq���gw��8zr���hR��}?q����{�e��p~��i��	p�eS*g��?o*�u(S�n*��Z�Ul�m��^Hi�񸑮Ա�[S����u�w�NW8�;��'��=r��W�a���;4�s-�t�ݸ磎�o�LÉ�� ��1ç�m�~��Ҹ���
Y*ˣ4�������_�����!���n�������ğ)߮>�+�5���OD����l���'��}p������N��I���)�����.��+�,�Ub�ZF��VW$��i.��X;�~�Szm�U����.�>]�i�o��ѡ�y����G��T���[+��i�'z��a�����<�!G(x��Ū�xG�k��*^X�&@_�$��Pt�0��8�{5�sR�ǟ$"ծC׸�(�53ڃ�B�^U�׸թ]~�r�G$i�)�'$A�z��e[��@��t�z��/Q�������v����h/�K�ߤm��ҀMX��瀾�?�N[9[K��/P�o�n�R�7��[��]� �-��K��cqzA�G}q"89�UG	�u�sTuu�wX�Ast'��h-0�o�Qs�5���4t/���-���r0zƖ/���ǲ��t׍��	c�FZ|�#;a+�Q���I�!p50��e���hX*ҡ�s�Xϛ�^��d����|=k��B̶I�;��ǥCِ�5C�����>ơ\�BԸˌY�:%�<_T�EF�h�x�&�94��J���Ɖw��u�<Z_�V�;��ķ�;�9�ʍ-Z���0�'���< 4�
��Ӝl~���_`�>M5�ۊΉD<�V}?��:~Ţ��i���J���(4F���a����5�VZ������V�i}h/���R(�yz������vd?��Y�����t��jRS�N��]DX��4��n�~����=O�*���C[��$�"����}R�d���) lK����(?waZ��4nͩ��K���������-���P2����:fC�(�\Q<d��~Ul�&܏x M��;o��A�AL��z�(ԱO;¨$�@d9��P>l�w��e�ａ:(���%v�'սD�OF���&���F�`�\:ۛZ������ۚAu٢W�����Z��b��n)�&�4q5:G>l�!1�e>>3�@L�M��q�@kq�@NU�9��q�
ݻ��T�΢�>Q� ,� D��	��k n�Ũ�àob# R?%-��[N�'��Ҥ���!�*�u��߃�Hz�1ʕ���r�2�{�|��l/���o,}�|�5ѪΙ�hz���g����ub1(��8v�#P�k�i�ʐ��{�xa� (�k���v�B��Jb.�����Ո*G�q幧C�x��n�&���=w:���kW�b��%�E��ɴ{Y�����K!�����cHg^�J<�yo�o���nY��+��
�$�'W�����£�� �?I�싶T�!AX=G�ۈ7mN������t�!9�6�"D6|�A˔��H "�(0܋�7~-Q�Vʿ&�����%�RV��J��5U���{�Q�m\��$�E�;��*����T�*��C�",����q����-w�Q�Q{2.[=��J�a�y$��v���)q�~�:S�T6u,�T���{�����+��2�W��D�`$�>ܹ��`�7?�����y�K.5��ࠔh���˵��,������_IW/Z���(��Me2��<�������Уڤ4E|A�eU*SQUi9�`��s��i�6qT����r}��̫�(�(B�~�܋�}��ԟxl$�8<o����}ښ��#7�73�n�/�ә%�H�}�МG��2T=� 26MQ63�[I8���ё4M�Q#-��D����L����*3��݄z�$m�v�W��v�mBS�FZ����>I����U\�j��Í�$}33CC\�1���H��������|��7���ER�m�y2�����Q2��� Eb�K(jE��hW�S�@�� >;~1����ĩJ��fd#��NG��� �x%��>D JF"�4���p��|��*�՟���A�p1m�I�J�r��pU��D�B�����?����m0ɹ���Ę!;��~G��k�v���8��1wFm :���f���!�����Q�T�I��U�H���{.��֦nk'��.0m��#�AO����y�0��С��}�gq�Y���vj�v����,��.!���+��E�r2�*�7y�F�ă�*{���G�����kZ��چ��7�9k��k`�>�]��K�
�s/���K��wA�/sX�6��>���(z�8�~]9g}�Q[#�$���oюNb���+�N9�0��Qf���������?�ӄtézu���-o3�Bn�3T�`̽�te�������=���\�&I�
G{����W�/��R״6�tV��O��O-�r#FU'4���*?O�5!�Ώ7�Y�(����pS��'z��̏�k1�p�ɑ�K�o���I3�������� 
gf��$<Wr��M�����49�$��	)�����~It�2��3�{�)�vB7@�7s��c��a}�j�}�ct}��4m�VgV4�C���_=M���qͿ0�L�=e�V�YN�ϫ¤%��`[F�A�0�g5}Vg�D�W�����,]���ųg�ߖ���}��gND����%}�3��"<�e�b80LUƮ��HsێȒ0A��B�0�@����Piᮻ�N�:zj���u� �� ��<f)��I���n�þa�r��0Q�6��%F+��o���ى���.��h:����?��e0��o�OjV�e��5��ǜ��)W��)~��LM�S�F>B`��������pj|���TE'�<I�%8�F����-.ŁrhtM�bD�k�Ku���2nV��u�� ''Ck'�j�z���,��"����EB�u���{t����,���,�5��cN;X���÷ӟ^6VU7���!���d��CX��c���?�����=���6	ak�x!.����-
����0M�9o8�#��"[c]�K
9�.C	[UV\��e��"x!W�:TF������l�9*/���D�$�4�*��BDmP��	ߠ#��S��N�;$��4nĨ��A7DIi���ش����G]'��-�B��a�m���K1� Lb�bB�xz�~�8R4K]��=�3ť�Y/*�0M�Q��'F�{c\o�zbِρ�qU�s\�Pw 6\6���ھEou���(�wbZ],ձ�SN��F�hY�f����sy��e#>E���y<���k��z^D�~]F��e4�Q���V���<�y
6�����k�V�l\(u<ޮ||�Ky|=FLڏ����1�GKk�q65П#�,?~G�Ԩ�#�Qb�P�)
ŹzJ�� C��Z��{�k���;��H�8�6�񾧉7w�  %� J�p(ŶV`��p|e(��8J�������y�X�k�������֛滜�܄�v]Bu�VEU���dЃ�	﾿I���@�i|� o��燲��5ӈ�J]Jי`��F�0���?�K�B��R�4E�� ��1��k҂���0R�b�2c�-��|:�.�g~*�Hs��S�N3F�V�|IF���%�D�F?�ix�4��ye>�X�8��&�(6�}l0��>mǂ��k��2��܌v���jdx�=F��������D�֯*�5��d�}<��8;���oG�����=z�
���6��?4&J|����a�!Xȿ�� )�6q�9�{S��u�Y/?3��E�/�q��ɭ�tt�����&��W�E����
�".�e�E�( I@T�����H�*A@�� 9JΌ�䠒��$�9����n���Ͻ�TW���SUӓq�+�0����@���Ը��o���෷-�|��-���vO���>�԰�T�%:��q
�q^AQ�=c�m�}�]s���7�#w_���	y~����
ާ^�q�B����x��]�@\�9L�03+�*��n�����Zh�uw��;��N5�f�J���'�9�]�|�Q���rT�ɦ5+���wY�^ �U�߿=J�k��rW����͝���K��v.��t_8�s&��u������P�.D�8�t����{�����OS�^���y��_���S��}��7����?�^9z5^�E���Dة�|׍�.Y˛�W
��++�.:��2��A�د�ةg��lվ�n2�H稍��&	Ҧ}�3�vg�u(m}�@�����Ř��N`���Fc������n�/�ݨ�A��,��z
STb�m~���ዛ��r�7k^�v'H]��ɂ7кn0ts�E���5�Ǖ�qu�Kۑ������,��l�Vwk򡬂6��4ӯ�o4B|�j��'�#��v�g�'�v�v�ۊ�)U�%"Dc%�d?���~�Fu�!Z'���Y�i��������}�+���%����ŝ��s�z���ʎ�����3fu�y3ЋjR�p��>�PM��mZ|�Ӓ~�G4��s��/}�XB\9��?�\�9��!�hy��gk��/p؇d_��]_��)�ZB�&���#Z�\�dZD�iKύ ���}0���T�E���Mk;D��D�_nw�������s��mY2�/<o<h��� �c0e<��h�M�FJ$�n}��h1�����(/x�i��!Fi�:�����l]%pcPDO�m�H���WH
��?X�.�����_�ig�����}kR�[�
�� /��y8��E��l��4+��w�M;�x#�f(wluaa�J�.�dbxn��4�����2z${%���������8q�����d�*����O�5���n�;�O_|�{|L(�X/��`(��b�ͪ��j{�T�L�'�1S��EE��Y�y���l7Jn�	��˭�k���OA�t(�>V�/SCS׈4�����q�7��,��B��6���I�Ш4�=���.+�T3��ZE�C��?Y6)t'FAL����uDf���W��R��=�S���M����tf �S�ЎsRV�SVR���C��A蒇M�%h�S�ZO|Q��í�e���'����@��p�ֱj���cb��ַ˭ϟl��2����h֗�;#-R��#���P���� H�e��1��ц����׭5�ow��	ʏ>w��u5�� �ho/9���ZJh35^�܏���+�)7]}���;��o����:��)h�M�c��d��h�Gtv�[��vT:��&�5�/��0�^td1{���N�f��)Q>��ҜMn����ֺJ�h�����8�W��x'cS�J)��J�v���eNA[- �4j��E���v�ւ���`'x����W��_�n�ܠU-0��Qc[���Ug���  �/H�tz9�G
�9]m�t�}��`U�뱐�~Ӻ*�f���.<;�`�������]d�X4u�=2$���2|�K`���J�;��9`_��VdZ�i�޷��J(f�nN%;H�&e���NaS����|�")�ՠƟ4��T�;X9<�u�O��R�u��/������Uϓ?_��:�p�Xp��[�W�^�acػ�X�]V��~1�o�5�y�����w�}�f��b�^����Ph�y��Ь��>;�^^f��ҫ緐�?
C���{];"Iɐ�xiQ3�8@�s���ûo��j�.x�m惥��y�}��:[=�CL��Or���8�,gz�%5����bp�!h�<������X�
kS%��V��<K�Y��c�u���;������O��]x����Cjw�+�K	�D���/�QA<��}X�Q`"���c^C��Ә���5U��3+g�G,���f<U��+rn뗔݃�МU򪕡s��^�v#,#J��׏#"�4��[#`L���+u}�f��$a�<�a��w��,a� �@ET4s�e���*@hj�
@h�M�O�l��zZC�)l�;�TӶ�^�,hz� ���㫡�j�=�^:��^*<{
������1�u] ��%�f�������op�X�7M����a�ir`����^�ʇgqm�w/n*��Y�!�N�6�d����d��@�2�!C�0R(�q��t�K@I��Ϛ��h!�n�r;1��b��	*�1E�������T��o[���A��ޠ��u���2��ܑ�����Z~�hH:^9º
3�u�,E��h^vO9R�Jn��c��?��o���H![����֛RGO�[��oJg�����oBG��>�ߨ��0�3x����k�xj�N{���r�@�-�aT�b[��r`�'���ٸ/�s H��oN:��kE *=�~dՑy
��x]Tp��gx��Gr-яo<��_,q�T�����,�V��7�%7^�ƶM�KknVAd�f��1(��l��~b�6L��C+&��c�	�j.b��7�!��|��)3J�@�T��d�LAJ<=�����Dd�T�w^^����󦼒K���g/<w4jS�$t����9ǘ���$�݀vZ]&ds�(�4���?\˅5��=t|�Y�3�5����u�qA�P�Q�6�~QH�30=������1���m��_r�ǟ6 *x����~�>ߓ�]0u��ZVa����IUN�+�U3�
�'?:F|||���sX�ΐ#٦�v	����p#$U89��r��a̙騅����2䲫`u�F�_�Aߒ����<�X����[Y�}P9�_iL�$3kDk�RH�A����>p/}�!
ȸ�&�΍�E������w�@>G��GVZ�Y{��V��ޥ���_�i��,�Q}ݧ+���44@Y=�۰�z�V��>�����k��##Ҧ*���}�v%Q��K�5�ZxM���������x ��wB��p�v��"z���
^dH�
��`j�t�v7T��'��甪��t;;m3�H�Q@�Ă�4Rm)�~�<&��?R���ӽU�� ��������a�P��o��4��Ӕ`Q;����c���8`�G	���@M7!����3 L	2̓V}�h�۬��V%��<���7ch)�e����8S�βֆ��
�Z��	1x����WW�� ��
Zz��\4Ҍu%t���.甼�K��Ѥ�/n0���(�^�N�2D~��M3�q��,y�)�c:n���F�6���eN� ��p�8-�I�-i=qWX�	
Z����z[�A�����r3��O��
`�c�a�\�~�h�C�2�/'�.�NX���9'V'+�K����.�v�X>!3�2j�dp8��`����B��P��,J���f
[Y�L#�ᢰ�`Xv"�:�c5 ��e����>��w�0Z��|ei�E�`O��qT���u��"_]�=ZM�.�ذ�2��\�`�^�ྎ�Gf���7��l�o�M4�� ȴi
�z	��t����|����ަ~�vWWCNtC�N[���{�U��	��[�
^��\���a���G��K�㟸�a�D��W��~���xo��@P�#�RQ�|R�#�n,g���0���\���ԬNl��,A�z�k�޽,-��,�/.��h|y�M*�
հ�a-�-�쓻`�^�,���;�8/WP���(As2�Aq+�[A���^��&�|� :��x�Ī�Gº��{e.�`�0�݂��z�A��<[��M�Z�`M�G�.XzGڊ>
�c�����K%�$Ô��vf/�����?�y������Ѿ���X9R1~Wx�j�p�M>�13����|��՗��Pv�K˪ǰ����j�ӈ�u�;'l�K+Ҷ����d)�$=Q��k�y �~S�a�_��"'*�m(|8�/�V+�l�������4C��h�7�Э�y������odےZfkA\����wH/t)����6��I=��vp� ���:P|;�0�.,�݉f�uXﺸ_�J���q�MgQ��i���:Пv����L�I�f�^�r��G�|f[X�w��n���H������D2��o�q���8j%�֤%63%=6�v�;���2����|�כ&��x�&�||n#&�K_(	��|�y�+��?��5"΢=F��?:�ef}�4s�ygvH�3p���|���h�Z�����s�?��N�z���QЪ��K0j�/����r��G�<f��]'iAւ_}�|×>GA�u�1h������/�U���V���H}�)���7����:��tƇ�$��n6��
����.C��cXtޅ
�f�H���h˚j�7Ո6纏��j2ɯ��j�T������3�V�ċ�U��#MP������֣�S��U��[��k[��P�8��V�Z�G��7t�E�ʗ>J�~�pd*x�CDT=�Ѳh>�����Bz[�D>7�ʇ���
y-���Ϩ�C�;�5����`G �c�`���A��������
W�B��6���=�Ǻj��S{瑭��폳��������D��#l'^$���*ϙ�1iAM�
:��3ɹ�S.�l!��V�W�� 'i��dD�w�*p}�c���Aj}�q�?���V!�!O�i�S���f��	���I�&{>0�g��U{������[v�aZ?��ƈg6��W$fN�H.����]�:�23M*hެz�#��ْ�V�G�����ں,4U��!W��s\��ô@sߟW7�����GV�=��m�t(OC~�D�i����"���c�G�VfI�$7*�g �UG����e �_���Hi�ɠX�P��=[7P�Z�&������:�� ��!�&~���'�F�j~�f���r-�3���g���<�Z!!��}v�ģ|����L�j�y$�T1V�i;P|��u�*<��-��-���<K6�J�֛u�hu�|`���
'��lפ� ��.�����K-��+;��IE�hN!��\��<�=m<������x�Bc�j��V��}HDi�ؑހ��7��3r+r�T�#�5Iw�Om�XY��!9�ܒ��L
��=� NQ�K��Ȫ�V��ֆ��.XM���Tz��.v��"�׿VL�e/���}<���qH���kH��`�g�]�d�����Ԧv�c/ë�֌�q*��{1o�`帖j���E�-s8�k���"��Ú�{�a��>������k}I3��aLe��k����������G��S���?��̤Tn�+n��l!��=t��(*M��'G��ۜ���|7%�"p�Rrm=������]����y�k�z��6/6�h�q�$|˒�]��v;.hk�os*�a�K(�	��oM��� �	}
^�w'U��̀�dA+�$f8?w?��%O\h/k��#�����Ҋ!�#[M�pX�6����&O�%̴�X�8���Y��ϵ��rM&PW���c�~�ȇ�:�A�`<L�=���P39F�qU𘛆�=�c[�0l�Cv�ap�_�$��H�����5�L��  H���"v��Y�V)b�xi%湺��x��d0t��Y0g��2��kcյQ@����Cߘ=�fa[�X���(�h>���%n��>*���:����Z9G��z�=;(vB��@��W�Bi��ʥ�R%
�;@VNU\�3��߭u|יdI.��6�6�h8솽���(�R�#��5Q�l5�y�w`�,�#��������s���X��c9x�Z����=�Ѻ�RG��m����SJB��aj�4��k�v��U�u�D���(���&����j��P��R��?X�	ܪ�@����N�w:��ܧV�������$�9�6#�Ɔc6@M��:5�q/�1A`Kq��>w`������!� UV��c�)��a���k@�C��&��U���!X�X'A��#h+dM�����|�����m� ��^+�V�yI~��
��ɲm�#�����S�M�*��Ӭ{�a'h�����{_!7[��3#�l�I�ؙ�A9Cq��[q٪�)}�8h�^�EIDHVV�;������췪NnXT��o��D�R��]�U��bG�#�z�&�C��|Pb�8�[��M�8@�ix���ۍ�݋��&Jpu��J��T�蘵S-����d�7es��N,��jK"?5��|\�!�
3�z���~��gL�P�EcP�>\!b��MYD��ph`n:���tN�w�,;4�����o9�k�S^�}\���E��l�[v�gE�oϚA�ʪ9��g~0[ëbF��]ѻ.���S+0}�Pn&�JF��� ���!�!�C+%�A=��k� `l�}�I�4{�T Z��}d��k-J����5{:,�#}�$E'y����Ǟ��/8��C$퍬����;n�>h٢(i�
�i|n K㐡�s@Tvjn��V;�qplG��áC��cIu��	�g��2��|����\>�$PG�-N4gQ���XD��<Ą���ʎ�Ab��%t��Y���h��YЀ����%v�ʹA���7����\��f�<���� `� VS	}Ֆ����~l<�b��ADD3v�j�j�V�� ��p�f��n{~됡Ҥ�̱��79\\���#�1���$E�xiS�v1��pͯ<�,�X�Wt�����HFQDM6�K*K�c�4�c��l� m�Ϛ������I+t�o��ʶ����܉��L/^�ݲ�=Q\��"H}&��E�+�Ӛ&H �M�;�]��UmĠ��9�����>�:��
�՟��$��|]J�o1RG"S���u���^��|��V�Vv鞙o��	NC]�0y�w|�^H	'-�q��C R�wE�՚���E䔠;k�&t�4xxw�������� ����Yv'~.O�#4��Z��<&J���j`�˖h<H&����R\�%�g�n/t̚��ȍ+��gy%I���@�H�|P��^�+FX�`<Ϧ���Pn���Hv�4 �W���h#̢�+˽4#aih�*R���ZU%j�&��w)A~�S��<�pw����A�#��+g˓$��3䠡@�g�{�&���'�j<6ж�2}Ը�����b�y/}�mh�ݡ�0��`�<6���Jjj��?L����)�!�%z?��^Q�������W�U�M�ʹt�3pޛ�S��̌�������0�,����_6�d~
��ϛ�d"G�C��x�����`���*��D��)d�����^n���c�0Q�Ȧk�;\�0�]g������u��̖����c�S�������`'�m�(�yi��լ���ÍY1�4�� �o�	��`�2#�Q�:��M���<�~A�)��/ESb��X�5s ��Kj�I'���s(��#��"k�%C{��PR�B��^ڌ-[����s��� Q���GG��+v�Vɇ'Gn�à�γ��ؐEf�����4��7��}k~3#�ަ�ޝ��}G������aG���OCV�)h{�;d�9Y��ڎD���y��5;�~�k�!�����t��`�KN��k��9fKT@%�ύ|����������86u�I��Gv�!Z�!9XjˮH=?����@E�����j�ƾ����|�=�`^�4eA
��BO��')ߋ�f`�pX��^�3�jy����5����$@��uy�K��j9iA(WqN��|���t|��CG.�Xvk�Ճ�b�Ƒ�w��x4�gl��Yt1-	��ٗ Y�i�*��%OU���߽�߫ۜ����E����p�L�c�%>�kdB��W<c��4�cu�Ҝ!:��e&⤫�CxVI�8E���T]+c��pXOJ�c�w.�)0j��6��4��
�'Dk+p�M����6���dp���F:=�
:qY�=Z��ԪuP�Z{�H��f-%�����fs���w҇��x��2O	����l�oq�i�^�G����C�!<wA�;�yX�Jn����)����p �����S �����=JH����P��jq_t�]+��\�nTv��,�@������O˭�9ORk�4$�,���4C�(���3���[���0�վ���H�r]2y�Z*����;�a5���T������ݞ�_����%z��`M�G7 �Wf�P����er��[�p�[@����_f�,7J�`vV:�����m��9#�W���/���YZ�+��������m2$2]V��W�'�vʗn'�ykKq��@�w\݁J��Ϗ�m�5���
d[A�w��piz5ʼ<���e	Ād�Q9�k�������γ�;ѳБ�᫢�Se���N�F��^�D6{�
�rǖ�L���OV��
nq��e��0Γm�G
Ι:�3�H�>�knrGO���WC�6	JƆm�\�F.	>ܑ�XJڙ��Wp�H[��_�>;3(��ݰ�CB��<�A�l@�76
�wǪ]]����A\Iok�Ƈ$ᆝ��?Y�t(�uS\�����\�	�Sn�'hb�M<������^K�uA�9�˚�R�ӿ��~*Qh������K
_Cy�B���Q����m2�.I��?���g��I���3~��y!����_�;��x*/�SՖ�z�n[}�y�#1"EC�i�Es#e��uh�F���-���.Jz;���p[��2|bk�(�^w�.J����v׊N���p�%�H���JՍ2�<�B�u��&�I}��5Re����hPb�X�N���Ty�Թ��#�[R9p�k-ēUFu�Ҽu1�T��i^l;X�����E�:�^T�.�P��։Iѡ\ޜkd�/�G�Ə���%�ts����?���Ks��m�\�xz����&����!aQ�^k8p�@ʨ�Nc2}�Nf�����u��|;�6Y��z�2��;d�v;[�"���Yі	��VK[���7)L�����D��ų�a��x;e6\�?�١����@��H � ��3e�͆I-���]��O�H&�MZ����V������/\�����ɍ'����o��́�~�����1S+���1�7g�K5�d������.!]�ߚ��}�k��Y��J:j�W����&���=x��\b�s[K��F#�6����;m�6ڳ�$)��й�X�#��Wp��f���t�\��	�yh�Q��e}�yv>uZ-Cw)����-\�n�q(�od[-/ufo �M��)������'���2���gsr�wN
_�^pKF^;�y���V[Y���~�y#=�/��k��Xg8�&a�Ŝ�?�K8����ĭ�և����<,��<���;u��1N�N�����s�E\�Z��>��Pi]3T	M�91�"h����Hd;�c4���>>C6���7�K0z~B1�U�R%-w����r��[�PUmE�Q�lC�MRg?�mt����{��\-�1vh1��[�Ha�?Ś�Ί�GG�.C�W�:jpH�#/_h��E���b}��_KM�ߤK�P�x�h��CB��\c�� �g�UrU)����e�8�ly�գ���Y�AU�����Uq�%+.��*몔t�+���rFx+ �1='1#"�6�!�/�#\>I�?ozģ�U�|Rv�YC��߬G�WXR�_���u�Hz�Z�
�X�h�{P5�U�ĦڈK��\�6f?�p��vp��u���{��8%��*-���~gi�J�m30f+@u��!���
W���u��ا�;�%�z�ǻuI�;
Ъ���xiJO�u�9b��]�a�òev!~�֥�ó[��*�Qy��j*�oe�밉��Yz,	�^�ͼ���߮l�`��<�5n��u0��q��r�XZٞp����~fmIF�/��^�n�y�*Y���El�)��,#O���ޜU�>��r_�{b?g�-�Q>́��6I����k�bu�F���*��ׅ�?�xW 6��ګ1��
N∢R��I��+���)Z��>?".Ñ*������G<C��{Ҹ*������%;K��IP��L>S̨�	�d� �a�/F��"�[�ӕٍT�2ˢ@�o?��%�u��c�^�񗞲�zOlĔ��[�|ccGh=�㧝bP2	�6�F\��)��>ҿ�M'Ҕ�2%��)��=����}�3�G&!�9f�]�a88;���-��B�������pp�:^�5Y0����v���aS�P�w�!��([p�Ύ��H[����w��8q8.5��?���S��X.�:�n��y��}��H�u4"�ɴŰ�bP�̠�J�^�[��)E�׉��`
���4�e�,�~;�M*��*�D��qO���5�!R����a��qeb�R�+���.%wq�g;!oiC�ۤ�6{GǠw �(�Y���f�~�������E=�p���c�m��ۈ���ד���9"�5c��Ha$���rpi��7\�x��t�ߞ�ۑ�V�s��6�6�b��k���;��N"�����L�$z�2E6KHwO���Zґ�j��N5��U:nq��z������la����U�K��!�rq��7�p���tS���Ti2��J7~�85U��H]N�'|Te����T��γ�r`Q(Os$G�����qi�LK{}��|����a�L-"�l�������������xڳ�fY9 :��Yv�f)�QB�F����+_�g�\�RP�
Иmh����CB2y���|�!Y�)��KQ̎7���Z���ZmzFN����k��}p��"�M����1�� ��T�C���/�!� K�ێ&�
��RWĕ���
f��{zEC�C��֨��j~�{�c��Mvވ�@�\̠��咰�*/��/��FE�lq
f���������ٖ�~YN�����WD�������jr��M38��j������?�e���z�"�
���cSƿ�r�3\J_����7x��
@�R)���A�9d��o��֝t��AiV@=H8^��/�Xf�(�tG��x�&�r~��8o�Ӆ������_E���'��;�}�i���MԖOM65Y�~2� O�\�84��u��sC�(d-R��gy	K/���~9#8M6	b%iP��)�����>��(8;��^d�T�UJ>E�;�[X����I`�W܊�0���3Q)��B�v����ld%z%�*�1�A�R�#�6�[T��:�0/[⃔m�qb1dMY�Y*��k���l���g�������v؄���Y��G�o5�h�+~L�G�'(��u�-��^=��B��"�R�Fl2i+�_
tts��:�s�y��1�?��o
�fgޚ�^��D:�4�˞`���p�뵃�KoM��60Ӈ�A3`�b��>�p����J.�+��Q�2���a�;�7��c�%"#kD8Y&R=T�#}��X1�$�nw��TI9�w��uM�-I��0;�4�B��.|+�Q�?dT`���Z��x�A�P�<p�3���F��1yr�1I9�Fr)��#0�N%t���_� ��J޲�!�B {A �r|��N[�kAA�� ��R..6�Lt�C$ �[;r�;�%M\�s�-PΙ��YS�%�+�0��'��s� �Hn��%�ft}��pȾ�����H���b*sSr��'�C�Zݻ'��0��l"ˏ/�|�eqW��8A^UlLh#���	���Jq���' ��+֐��m������Wl�HJD�+۲�TZ{ܨjS��5��h)�88���V1�?��B���'~���ɍA1hpV0���S�ho`;ڈ\��'^b7A�΅���M1���^���,��J��%D1C��*�g��/q�NN:M2zQc5�r�`�<��=�'_
��SX$p"�7�#	f#��(Ys����#Fp�6��:���5��M���
�3|_��W�S�1���BSн�;��+	+-�Hz�}�*�8?y�Q玖3����R�5Cyi�D��!���ն�Z��Ԟ���{�Z#�dq�u �����Ր������<��� �o�R�>RJI����+��i�E��d��V�4�m�����o!�7�"�ر��ˎ��+T�|K���H7�V9�k�%�:!�v^�����xQ��XŌ��\m�d��*�,������}�?������V����-4��	0�U�H\�.#�S&cn�@�v{v�o��)�S��s��k���B����m�=�\QG������W�il*F3���� 6F���xh�Qe��l���ь8�HJΙ�I�s�"�ܐՅ�߳�w�fX�?�ͥ3�c9K��ݚ_�ڙ�p��A(���qA�d�=2�rC��[�%6+��'��h�2�'����Cs�ĸ7�N+D�
��h�Zm���O ��F�˕�b�5m�7�ۏ~���Z�߈���.�x�x]Z��S�Қ[Te.����(RR	i{������aɪ6�Nd�E)i�R�&�VP<n�wd�:�����4g��{��{l�ς-b�u�_�\��R���r�֤2�$�")'�Fpoρ�]�͕CU�y*�b6Iˌ(�޲�Z;#�+�[i��K��|���X�e}���%/U�@ 9._�N�cWS�b������aA lsѩ�����Ǔ���xࢎy*���.{��	���!�m׺��nP�����Fy��+3��3d���Fmr��xz��yz�x�9ϖ�q.:�q����O	 {�?"h��f�����V{�V�0��S��~Do�?�>��pf�yF_��ףM�(g]X��P� ��2��%uZ��=�Uu��n�-�=?��'�\T�1�a#��sM>��6H�z-�>�ͿG���P�tw.YbӘ����T�9:�^)eRO�{8��~�y?4H�E��WX����VV��A��Ε�'�����=C6�F��
� �d�j����]%�~��-�1�������#èE]����Z�q��q[_��v�����SKM�Pm�5�zZ�j�����Sv�F���9U?��a=B�o��g��!ݺGzWg�� (�SM{u��k~��&s�bu ��OA�ow'���욭7J鼦��m@�J��>bM;�����8%��؏�h����*�X�8�j��T�uR`�bu�G/L}`��|~�S��R&��г7y�ܡ@��(��0w�[��%��Ɵ��vf$jH�b�%'�,2�W$��44_R�CFԉ��|n�Vy�@Z��
~ъt5�֜#�d@�{ŵ,�
��4�8hqX�OTv�q�rƟc|��W�HCU�h��'���Z�Ј�AQ3-�����~��wF6Ih�QB�O���Z5.W�J�eKOUq���%�)oT�pB��*�pŕ��,�8h�/��	��=b�j#�"Qn��;)п��Z��~�\��Q�K�n�U�L�A	�R�
�:��!B�>t�ދ�.A�7��ȫ%���8.p�`
�{�4B��{�5Z��3dּpń��L-�.2x�P�S���q���f��_S�iځأ�v �A�h�@�bhm�Ju��������w�E�pE8_��^����%JP@�[i�k��~"A"A�eǞ	���H��.F�n��b+��#�� s�ˇ��ࠐ�W)&}��z�Ҍ��Ҏ�a����!3��d�؛#�oP@�$��:wc��ܦ�:����Q���!PTP�lT��"�?��݉*��m����"�n��0q�M��c�ه~ȡ?�h��⦾�8�m�p��UX+��S�?������"m��t�6��{��Y�_�=�̮ߜst��P�!^�x��L���;U���������1GȓB J�*r�ða�ӯ'�SU����P�l�C�6Q:����� E+?��b�6T�+Hͧ�f*�MڠyAjEE�E ��UAE~o����㭠�g�>hb豓��]�	S�� ������N#"�:�����3�V���et������'��d"L)�TJ�NB������j73���
㻑��	�B�/����1��~0ⱽ�-�#ѽ& �s%�r�B_@�����?��,˂��V������BۜȐ���	i����gU��ʵ��؈�h@�x�����7ȯk�ǡ�
��z��_���1��՝���u����+$hU)f���|n;2mY����[`�]L3�@�?mU�%�C|4 |,��S�k��Q�l�U�NP��E����P���z������Ϭ:,{��C��F��o�H�e�0��T�D��&���q�@��T��#��Nn��� ���%�h����OW�I����~�#�W.�Ӄ�q0�GDƜ�R�8�#Ÿ���+te<peɽ�1|�g�j�,C�/��6���G^2Wl?�����ϡ�X�W����h�kw��u	�{���%w���M3R�
9�9����;�V�L���+C6����g������/�5�SCB@���\��,�|`UƔ%(г-o+bl����L��O� S����=��6��`�jëeK|*��l�D�u�{9�0Z!V��ݲi8���T���	*� ���͉� ^fZ0B����ʅ�	Ј}��2�;��-�Bn��lu� G�V�.�E�j�"���ƕ��L|U�t�_ѥ.�̰�*:��[P��m�E��ĖĈ������V/@�7�#ı��̃X�8/��#�nhN%ץ�dl)~�05�f�g@��j�	�����!\�ʎ��.vk�"M ��JH>O�}b�y�"��������!!�eT�>����L��x�i��3a���X]_[om����uE�� ��j�2��B\Va����P$ >�`P�O�����3�g��fsCTڗ��!f7m��H�?��ߵ��G߹��R��B7���_-�?1(��Ȑ�3�`ۊ����m+��e- 0��π5�by��<	b�����ܣ�Ou-��~��|/�MY����F�B�!��Ȉ[S4l�h�h�a�y[SS5F ��[m��-67� ������x������ݣ4S��.2S��qP6<f���o؀.�(`���4h�޳ 1�ԭ/X�G��z�k̍��Z#`��F8�;e�S���%Q�Z�rK'���- ��Zܙ��,QE���Y��W���aN��{��
�`p�̻�KU�^@�@U��mc�����ݿ�gj�e1��� ]� ��:U����.\eW����s�<u�t��4N�Ha\���*�KY�*sw�4J�#�e���=��3�����?�Z��(���ݧ���$)���9D�%���yt�N����W��=Q�dd.n[�t�p�V-�Xu��>�S������-n�!���x,�m�Q����Q�"tC���) ������)��h��[\:�wu��1\8:J��}���=�y3����I�0Zu0[��8|�G�$Ֆ��5W�B��bj%ܺtXMH��S����m/�*����YhMk�KO�����pe�[S4��zB]&�O3i�,��Ok�����4aM�x�#��`�����
<76;����p��K�U&f��\M�"U�|��з����;ɸ���+����X3�ʣ���1K7q4�~pE�є!���U�A�-Γ1iD��cm���h>J��=	.�l�b��*~��˃&ߩZ>UmÎ���%Or9%������*�����_�D��CK�A-����U����!��f��aL����˽O�UA�z8�&�P���ϯpd�Î}N��(`C1b���p10\�;�u�9���?#7�����2���a�RD�\�(�ވ3��y�c&>�Sz�p��O�V����n�8�ޤN�"�
��B�Xe�'Ǚ�3� j�j%kw�/�v��G�\�(�aI�����u�XE]n.j��Q<OW�\�˥�b�������P���a�����أ����mQ��ә��ع��#;��l�LN�]�)��ZΡ��ǿw61�|,U����1$컦B��ッ�s}V����&ͤY�FN<@���o�Rp�Y3h���	/ٚF��@<)�т���D�0��&+��χ����aW"V���+Ή?w����c{'K��L�����B���H	[�t�$�t�D	pm�8�%��]�߮��+W��mo���M��8�SZt�3���̠Fd
���?��Ҷ��S�ԣ��<��"BHHН=12J��.��V3�Y�n���?`�$�s�{n�y׻%�Oc�)>�*�<�\���~�!�p���w�z-���Y�~��=mf�p��ċ�ʏ;\���_:��"&�5l�i�9�A��(-X�e�He�$α������2h,�U�nʸ���(󨇥�>��5�0g�ܿ&���C:/nW,��W��5�ehЯ�C���3���t�����x҉���0�f�a]g�ց� �0��G������X�����Iyx}���Y{s̔�����犻�pX7r�'�aU^�Ē�������UM9�((���e�II��U�>�o�/���
h~�<��񳦮���7̷�$I����eУ�Z�-�'P�$`��0=���a-��q����3�G �Β�]~Wyi���x���4��X����1��JSH�4�(�f{$f���'���E�Hm. �����p@�i��?*�#�Uq��\8e�xo�����ar�$�K�G��p�h���]I{1v��T��XA�'h׊�ēE���6:��8�H�j�����"��4[]�	��Ұ����Ui]�q3`a��j����@��̞����[��N2 �'���˞���\('�O�"�����~=��>f7���>�`���pS1&c���ՕÕL�-d���Z�^���E�3��w:I;ے�]0�@�7�+�N�
�;r�@c`n�޷�Ѭ�;[�n���v4���_qÈ2��7�]$��e��t+OIZC�A�@�oE���N~��
�pқ�	gpK#.�&[��C�*Vop8�x�P�@��e
���g6�oe�3	�G�����s�hV�t��/aO����p�E��+s~��ľ���\�~�����S'�mVlk��� L����̹��wml)�ZF�I�����!ʶ�#��?�2Z����/
�w�||j;ȉ����'��].!�_]���-~��$�ϴ�I�Ǹ8�?��ߐݐ!G����̴M6}����RQ+ �|�d��/�K�-l���Yo��'�z�w�3:�a�ޜ���2�˖�������P��Ԕ��l�;��T��	�.���F��,i��xY�Ld��S� �}����J�-5��;����Ko�%��U}_#�����'�fm!�ds�K�P�}�b)A��g4�^�)Hvs9�MZ+�0�����p�*�����B����~�X�[�;e��ʡ��G��#`�8�5��AyIz�x�YIj11��`�֋���eYt��RWU9��I��/�@�pX�$������J�|P]=��?�6߽A���P"���G��ey�	,W�= R8F~���� ��y������Ǟ2"f��m�X�#F�ڽ��Q�ꣴ��[(�vݩ3�1��nc�Kzv�$1e�( �a�X�w�2�^��\��$s_�g^胢֐�~"ހ�S����aW�
y+� |]���%{T���h_x��x'��{�¡���a�/���{N�����c-�{	S��yW|`����$�)����5��`��<�f��}y�/NEU�]!G��3�~qF�D�h��O&�#��i�	���Ͷ"%C� .��4��{Z�pC��o�����k��� ;8
!(�;s}�&s�����a���S	r/]�Q�j��4M]]|��XT�?\�o]ue����؀>���JY���� ��"���PЮvi*�a�=�_�L��>�#bI��Q'
�,�|�yB������PQ��s��#�+E����*fM�d媚��tS�<��HH.������Ćy��$~ڸ	J*����Pƿ�2�̽�q7N���\~E^ޭVe����% �\bt�@R�]�,qϻ��i����a������a2�5� Rd�(Z���Zx�b�p�>��m���7I���C�����\��p[�$�@�����&g`���x֤��0�ܭ�	Q��̮��cS7hQ[������K_(ퟱ�$ƈ{|n?�$�M�;���	& �d��\c��_�>����\?�;#~�f��	�e 0YwT�^�ۗLCxn!A��#�3s����O֝�#F��2�M�>���ajʽ'���,; �e��-�}z\�,'.�ZPlh�~P��bx�. �oS��m�R����A���L'CrD�t"���{E�����R�s<�Mxp�����Ed�!���������D��蝵���$�5e?�g\}������"�/�H�,P�:9�{n�w�_Xu{��#q�,����<�����u�P����ఆ?s�p�/	��Xº�Q��ѩ�IG��編�\`��}fh�E��/A�"DV'�Y!ｭ�
yt�@<+���D[�qcd�'�"�I�n	9��oV��W�ЗJ�}��@��2s����l�G�i.�笓xW@�`�vc�}�biU|�K�/N ��j�����>Z:�����?�PI��:B�*�<��M�؇�'��,~>/�����
������&��<�٬Q�ܭ7�%h
�u·od�� +:�̋
a���,j �'B�{�ϑ��BQ,����v)�� � �^ �~��lİ���Vf��-J~A����L]u@T��vX0 �DRR�t¡$�K�Nghp�I���J�J9JI+ �R�1���	�?��}���|���n����Rʺ�B���a]`d�9W�l�9����-�qr��DQG���_~�oXx��(c��%ٗ,BӢ�vP�� �/�f�a�#��h=���#>7�|�>�l�/D���{KvP����L
�RI��[d���bo���U�D~e.��Zwy؞�{�A�����;H�H:N�؝� ��-Y��62Ia��Qu���ٜ�t'�)�	���S?Q/b<���T��WV`����_�L�U�m�r�4�˕ %��<<3֩�K�w+g�s�Q�?A~
�~j��؂��&!X��.n̘��ӿ�X�9q�m�� 	������Q�W6�l�H����w��jNk�QO�h�PXe(B���/V��B����P&���Ax���{�*(������s���������!g`�S��q��s���%1¯'�	a_,8�Hm����"4�Y߷-m;/�����R�������C��y.�D���Y�?�E����P�؂����|*2g~j�2b����)�P�m[�t�0DFE�';a�����U00���o�9�a�M\�YS�&�-�C���Dq^~�/�vp��!%䍬����C(#ť��3C5@c�;������KDo�,9��%�_����Im�E �/�1%��-W���|�a����vh��~y\�U,���|�k�E��ge�R�D�Ll�;�5�j��֭�>��0��-�����:}?!]�X����e���6� �Oӌ���+�?3���C�ߞ��S��3�J`�z��D���z�?�L�L/��-�$��^͌[�/��c0�Y�U	f�	�/��o��bo;/o(���D��+�Fj�OR��0����c��*?��f����� �Q9b�\�C1��l��wz�f4���!0�QN�j*�:�s���"̤��S헛SR:��9��}Z�&��bA�i�$��m�W�4��q�VޡKꖗ@�]�F����������Ì�N	X�w��cCܠ���τk:��8�5TTOgf21n*]
��7��6��V9�BUM_�t��kG���>��RX9�8�Q�Usv���[�Ч8s��i0���A�:�~��߲��B<�[�g�Ys�O!W�Z�� !�/�
)P��A\C.mO���fec�3�ÿ$��2����Rj1�&�u<� ���R�&��	3�iĖ*��p�� M.��)K{����ɴ�M��p�?L������+On�����ު
���t�;�A>wД����"�@�/'W��*�����h$�{؟V���$�gc�~������"�Tf��b6�|�,��@�'y�����V�+8�u`�C`߃0O8Y2,�U��"`����ŗ�>_֍�Dt?
$��v�"�/��oA��&
f_�8��H<�ޝ�fq��j���U`��F_�Z�i־T5����wP�S���/�O��ւ��a�~�1�R�����˺^��=�կs9$#r��_�@t�W3n�J��̏�����g__8��t��{~&&��"ࣗ��O��6�)W?�P��\���G���G�ɑ;��
��?n�ɱ��p֛(J~so�S��vn�9�
8��!'��!=�Hz�*B�n�jt�*pΏ�'Y�9a*)A�o��u	oPoh�a���"��KT�;�x�=v� ���X����9�cf͌,5$�������K���/~�O�SL�|��]�	��	O�[_�xs��\37�(hH��܁�vv�@�����p���W���7 ��9"����FO�Tn^�[�m���~���N���'�,.Uq�1v���u���;M�Ф7�l8�ʨi���A���7`!q6G2�%�4G�6qW�m����~���R@$�=ZZ�Դ_�Z�<�.鸀� 
L�y8vX1����<q���Nz#羏��da&)�~�&��O���{.}l	�WaFP	��p������iPM��C%�O`�p���n_�[Ҍ�$x|��Y�uj��bm���ė:&��g� ty=$<��S�LlnB^��&2��Oc3��������t�_�]H�D`0QY���gc��ܺ���́� �X����$8l;C���@3����
Ǻ���Ӽ�4~�ơ1*%W��YR� S�������3e�����4B���o-�O5���
R�.9^	���5N	��M�~���WYW��|��c0V̚vi���$v���#�M|��Lv���7�X'ر�ڂ��s- @��]��~F��N4���W���0�IY|`���O�m� ɾ��\`�M�`l ���`G
�[u��+�B3�q͌ǥ�g�r{���EL9�&���K�F�rr?+mKmC�(�OgKjAH�\�5�>�D���$NJ��]3
�6i�6�mA4.ǟOs�q�&*��ۀ<^q�>�yJ �;ks�b7Wx�p�� ��/�М0@��@���$%t����uzv��7<�R_(�+��H�Rf{2(x#�b]�rNKJq��W�D��a~����]+��!�Rc��\��}��`��X��b�Y50ޠl�D\��b�#��%6�|~�W�W�P�^
:�� (K���������_4��ȬK]�řH�1�1ߛ�<3:~:S���!^p�e���1�6��r�b�?��$�ucB�d#	��Ƴ��1�3��fu>���D"���wnճA>�d�d7(r��y��e���ݏ��Zy�oH����*�Siߐ_f�T�����?{Fw��D�,;�]Rm,E ����b�O�ϕ�,m	nঌ� �sx86�{� ���#.�-=ҩ�о�I�+��aﺤ�k{�����@�c���fu�a�?��P�en����jOpM��=���A&���m�I	@�a2������Wx�_�������`����g��	�U�_�IQ����,��P�'���r] ~��#!�։��[E��dn�?��IP�����_�����J15�ҳ}�OP�1��_�fr!J� a�Oi��ro�R�8|���y�O�&�������j���l�!����3��G��U���w�M#@�	���m�L�O=���)Yۜe�Hztu"-��>Ōq�m�)t�K�t 9�֖~�Õ�4���.7Y��)�Z�2�><�wm�v� �i蚍�7_m_XW��U|\Nx���9A��2�}�f��)$��?���X!���G|��������ng٠%�<�[���W�V�ߑ��^��)6�}�L[��
yYy���`6����"�[��
ӛ���O��5R��P� =�Dr�|��'6e��,߰�?�<�ݲ�~C�=+�N���_
��Z1#̓���_���(��.�Cϱ�^S:����G�Խ}8�q�-���!2(hq�̄�y���qi�@�S�Di���`����߿�x�K�p�8��}����OϿ�L�ކpp�i��2
ZR�]=zUwh�nnM��;Es/һ�4�
ή��p!>�䗻��"���w���R�,�A����~��i��No����S^�Z+f��I�C
�qT֘^^9���*�t	`[; '��s�g�hx��,u8t�9�0u���_���=p�}Ph��`����d�Z�jY]H\XuR�da�����#�u���ƥХ���������BЍO�����E�K�ߗY{���`���[G����eZe��S��%���y�-���&�,���ss�=��gC�!�ҭ�j��8�H��g����F�9�R��و�i	�<��g��h��oIIP~h]�B")�����b���1���I�b����s�}�2��b<��IV�;MBc��.��)s��с�\=S���b����́m;�)���'����u�������Z�c�I6�!1b�Z鶲��H$�J�ѯ�cV�eĶ��S�r`da#���-�v��$0��Xr�W�N��NIf.�:�̼�Xd����!{^��V.y{��6O|T �;��l^�,e��]g��1������n���y�����|��C���	�W��W�9�����U�b�����p��
����d���Њ��Ί"b��G�pq������n�3%�D��zMI�
cZ�H\�$��Չ��b��EͨS�	��5BYZ�Z�*u��U���2��ᴕ	���O{�i�S�h)�p0sCG�����𩍚q�9l�%C9�&n|sd�_��$�:+ځ�eo�D|I\JQe�&7|�Z��t�0	���0y��і�.� �=�}���LY�/xx�����{�A��Uj�\:5�w�V:(�x�LW���|�7�-d���{�/�Pu���$��6�b��b.d�C�ӣnb�U����}%�*�5���[�0Ã{��b��,޲�v~:`��a]��W�J�Kѵ-�0/ר>c=�a�(e��%���qӵ7�|���O�F/F���_A��L����P�ְ����XSM��13.�,��kJ�X�=�^�Ǵ�u��`]+�N�U��\5��{Ey�,n�=w<?�E2���JK��},{��;XW���xW�����x�����Ɔ��"���v8�,�^�(�ޅ�Α)٫V��tt�V���y]>�Ar$T�$l���V=�i�����1�|C,٩3^�������V彩X�0탦����?/E�GWs����v����+ޮ�t}P������a'n� �g�z��WPH�)G���ٯ\�c������ԧ��M�#�m�B�{{�Ge"����V&��\v��6n�H2�[TZk\;��Fd��G��祐���_y���,�Y0�M{{�k&���/N�,���Okq�۩u�q�����G_
V��$1fKu�J�4�˝9����QE-o���d�, ����
��OW�/7aQn7e��O=�ն}{'(HmQ"-�`����9�Y�H⛀m٥d��Ecg�l{����Cn���˸�a��'�.րxt���� ����3BB���h�w�VHa~��YD67�F�~:���}�Q���ۂ�#"�Lqsz����������Ci�����տY�;y����-��H[I��J��N�	��&����5�c;�S�ʝ&�C�d~N��҉M��C]���z����F��0yb�i����H���s��fZ�'��1ہ�����˔��[e'h8k������z2N�(?��!��`���<�Q�MS{���[���e]��o!3��I�����c7�!��G;.�� �*�������o�MzN���2筱ԇJ�2|-�<4v+���󟌚Ǔ�ͣ�<;���'+O/ϔ0�!_H�~̶�j��n�"��6�<,��J�L Ǯ�p��V�z�D*,`FeZu� *��F~���X�I1}9y���Q�D.�V�v3���zdb�i�����f��Aj���bw�H%������.A�1��ei�.�N�Z��/�6�4aI�`/�fwV6X졬	f�ae�"�6fJ�dE�dV%�o�;v��o����e�6��n�0�̠s�IVo#��N�z����V�mm�33ҥ���^�ܕYv�ϝ;�4hB|,��o�`�#��♙i+��*[��1���s���xo�9�%�{��5
sα�h�;�Egp�[?`� |�1��|}�HJ���?���w�J5<D��:���,�����2|2�� ҾQ�$}���H}oޖO���AP��%V�Ud[)���ze�S��?k��p��=t@էp���p�>b����	��9[�؇��o\��H�(L��}�d݊��o�#�!�sc�s�����i���r��~��%�%�4eK5�z��y�EV�k<%��P�]�k�>ǧ��3�% ��� ����Ǚc��Ŷ
�	��z��M����3�� ���D���n���\)p?0\���b"���:j�_�����v7j����?5����#6k����N�z��������Ԑ�<��8
}�q{�sdax�5�^���U����jքӊaoV��Ɓ��|�<:F}=*E��=$��2�Ԓ2U��&�߱��)�$�]�I��o�A�<u�x"}�}�Q\��BtEjz�`Q�����=�օ�<���VX���w@U&�V�љ<�
��-K�ו]��؛��c�׈�;I��~0��'�z�7����B\�eҾ����Atc����S���祈��f(����u�=�1��������j.�5�}*��p��@��7��2/�o�܇t��IVla,���>��9	�w�7���|�T[mqAEk��`�T9� �%�4�X�S��\�1=�����1�@�Ȣw�T$��b;�����ň��Q>�����z5����}�����jJua"1�)9a��<��CS)S|��6��N�՚�AK��MG�d��er���|�}�e9z�ক��7��߹/$5HND*�j�I�l�Y�
��o�/S�b�^-���⸎:oU�h8�K!�|�1j���>��)��U
;��|�nm$����̣�+��*`��3����u�*m��D>�z�;�bcm������#'��u��aoR�L�M�w�/���t�}�Ƶ�݇��2�m��y�ɝ=��H�mjߍ�t)(��{|�v.�$�s��h�R����D��,�l�X��yO
�T��~�A�U��X<M���v�/W���5@�+u�
*H�@�F��U��:���P�}�t�0e�u�������o�Bg���7nSK��!� N�*O�m���I�f� 3-����5F�a�J��)�=�����񙙷�70��F�}�k�����у�E�����X�_�OO����-Ҷ��${�<0�����s� M{{�����|�T-������"?���)=��/h�kKm�S���q���n�O�طy�,9�u���d^�Ǔǃ<�\��d��9c[I�j�J�El�i������#P0�@���DRC$@�@�v�o�U��Bt��M��Ӕ��)�*՗�MK`(�6~��$Hċ9FU���A�j�Ȗ����� ��C��6y�6]��qn�N8�Z�u�fv&jɿM��V���ci*��ذ{��ٰ���M�t�I�����KΫx.��`�F����Wcp6@6%����@8�DӢ�@���?t����xO{쀿:���-���?�ȜE�������$���������J+b�F�p�8V�34UWw�c���sD��̰���� ��~/�t�+O����M�\�v�^P��]�R(���G��a�64�(n��"��t�A���$&���̹J凗���n��sq~�p�L6��8l��K�����Rڹ��2tԽ{"���V�5�y�PG] p��%P��*�]��_�tyvb%e�l2,�4�nz�J�H�����O�Ɂ�y���BS�lt{���{�W
�#�()�=B��!����k��7�	� ��϶���a^�ߓ��:��!���`[�k�o���'�㊵LÞh�j���
_u�f�	�fF����"��!dB_��X�m��M��>�i�ݲ&l�1�^�I�X}�2�2%��U:r�����'w�om}n�z��D��;�e�M��U@@s _d����͏+)�wJv������3�i� S����,�͖)��5�{��\b��*(��Sv�@��&���%�ߕ."@�.9�4.� ����I��TS�7f�v��&��xp�7��w�!�5L���Y6�O� ^��/tH]��ur�q��0ff�"�f��n��h��.x��W/�����I�>]H�TM�Z�IZ������O��nMD�8��n��K#���(w��� ��t�z�|� ���ľ��U��/m�;P�=��_���|���2�w��b���+�i�v_L���'<V��9������]�!��x��n��T�5��l�G�z��c�_���y�w�������|�}�,��!���F�L?}l��;��=c���Q��LS��W���^2�6'�M\�F(�t3A���\Վƀ?|�S���p͈D�����lI$��_������ܞ�ʌ�ݮ�#�b2�ko��{��I�қ��E��Cc�'s��n�m��`��C���I{��[r$؆g���΍Nik*f�Pg�2�g\�Ūu�x��2Ew��֎�������wԟ��V����5���nh�U���ů����ly9i�����[[&is_�g�*Wn�)��ˑ��Y��8o�g��:��Ԫ������7	=��-������f��8�����i�g���#�ә��E��F'��^~��d� 3���D�(�WTaBf-���;t�+;�x�V?Ih�����AsL�s��ڥ�/��YF^ޛ�&E�2��`��#�ڣ�o�2� �0nԔ]�U�9���k9F5�^ǚ��6[V�
�fU#�-ON_#��thY��P�EB�S�J�����dN�J�ч���=����"���Z����R���2���a�<����'��$:����bA1F+Wu��n��h;_M?�>�u%�����/ q�U��Yr�%�r��OZwȐ�#2_��C�4�3�F�[ /��E���{�wW�����F�Kx'y*�^�;sn� ]v즶\�go�	�+z�٥k���`=����_���!��N�S��{��/&�����[oR�z�.g�t��mp,���*ն��$=aA�i�wz�p�ra}G�p+=�r�V�;��V�8s��%�Ǜ��d� aS}W��m]���d�1g�;-�s��n����rH������n�PHt���`���['�nW<p����8R3A�������������4]��[i<g���T�����w�3����[11�d�}��mϒ����=5cg�2�g��*/7��$v)���"�B8\�b�+�txl�H�\�j��^�j*�]�h��eC.�� �2�Or!���f_�\�"�h�r�?Xa�����i�]�X��\/9 ���3��,
��R�<v"���a��kJ�x�&��5�UT�
ǹ��9�cQ�dݥ2��D�K��	�h�d�;���	^��KVk��>����hIx#�a:����)�m7��{-��+m!u���c�Au�		���,Nɪ�@J�`s�y9�g[��lV:�H���qj7��#���,6i��w/�*�1oU���缑�?H����x�& uK�ɗj�+?�Qƫ���=�V`�]-´N�K`�����p�6Z������	�PD��D�Z���d#-���c��eco���hM U�𬻊G�c!"B��=�_`i����xH�X���^.i:��2����*C~D�F��MO[��3@z��I������kݬ�������Y�t�>)�
ͳ����t��U�YVȭ���ο��O�>�ok�ǟ����S}U$}���`f\��s���"���[��^�8�Œ��%���eKN��l����"8�V}��Z�14e�K6���"�i&��E�<�	�6;%X&(�/Ye�4��th�P�����µ"Y��DI�p���������=z���g=n���刴hgo�5���K���9�[�9�-s��Y��P�~��"S[��cN�kI}��	R�)gU_��,^xlw^	t�T��;��_3꛳{$��:@ċ��r�{����mz6}];�6���#���5ԈW�7���4H��D'�A�=��~��&��M�T��l�4�/�~����T**�~{Xd�!�z���MR�h�k��\���	ګK�ު��*,�/b��(��'�.�b�Uz�����l�	Z���;�=U��`[?`�]8$�u�}����Bz�9��
;����})O�C�]5���5�1u7n�+�;No���>��tb떣̿��C�V�S?��6���q�Ր�� ���}r���Mኼ'q����yЄ�.��n<�6�?~,WcI���a|t��xw�]<i�Tl�(.�	4:�@�`w�v���p��=��m�r����O|��k�1>�����ȁd±E����i��@�Z��HU�ܲw�D�swγ�0�'/�uו0���s1�ʌ�>?�[m�,���	�jeM��wT��$-�G뮪×ɏq�o�
}~���0_�]���;[Kw~��V�N����%�Ծ�O'���v�d5�����R��l7'�E7�?�z�M�wG�N�В��ho���0���5�x�e����΁]c��EHºɛ�k�	���Yp��o�I�����6��ͼr2I�#�D{e�ޖr:�j�B蜜�N�i�#{��o�:���v�q� ���y������|�`W磴�U�%�?6�.���WR���C37�����sA{\@�lmR�@´+�a�?��0oVDk��.P�\�[M=K�hY����xix��y�H�R�h��s�>x�LI�f���Q�V�;h��J,@Ih��בx2�.�9JJ�j����?��G�~��2蟲y�<%�䔅/	��am��!����S��c�U�w�n�.p�\8D4�G���k�� ?������*e&�e7���_�Hz�����b�\+V�.��=UE���(������c������X�;�L�^7�|E�X�i�6���8Qf;t2(�[�T�2%2��(��w>|:ڞ��]5xZ@�� I��X-��T�����R�Ʉr���gLg���|��BW�ܪ���cP��	m��'I^y���bP&K@�t0��:����Xh�����F��ٌX�p>9�q��c�j�j�_Kŧ�u�����Kz��f�{M���'9�b���̹b�2Z'��3�:��I)�,����cE�0�-�:	.'b�`$�ѺqiZ��	\tZ{�0�r��,��Y	�+K!ǂ��L��V�%#���(§|��eo�sV�����������3��[����5���br��c����Hi4`�ד��!Z�K�%<���E�Zc=:9���}�h�c��	�l� gv��Y�e���6��-3����'���bRg8VE:���az)�����i*���z�1�:~B�)���N�6��,�i����iOc��Ͼ��E�]�w��X �qy���R:q�� k��f�0�ܣ��Xsϔ	�n�}1�����a����K���� �.K�tզ��v�۪��3dŤiK�a��ǥ%����a�5����k� 9����0�p�[L���-	@��O���2�)��1rG��a� ҂��~��
�U�'���un9B�%I��٠^K��6���÷:�	7ϖ��:�u���o<��nV��ô6k�)V>�i%�?�m�W҈�V]��ꔘu|��B'z���s�D�en�q'D�Bn���83�_���z�,��S��=�������s��sb)�M�*�x�)�E>a;�?����NU@0}&}d��.���S|�kί��
�5=�"!rv����j�<7#��x�#�D�o����7�ky��y~����rm�����x�|:R��?��Oe~r�� �I"%�2���Nx4�ѥ6DDFz��I�\����ܜg.qK!�
��3���lМ�t
���(����p��}�qbz��W��-ۛ�C���W(^t7�a%ÒW��@uC� �jo��ѐBB��4f�ƽ�����#����v�#��w�,L�֠q�{���	8AB�&�G�kl8LT���Jp�O �x�\U?�*/bK-ʪ���cD�G�|�{2����:� ��s.^�ȏ������	��m��J��*�!�S5{\7<,���zb�;<��<�0L�� ���?u�ܼ<�G��W� ��FD�8)U[��h@����۳�_v���/� T�./�$�h �z����#�?�P.�_M��]�#M�2dq�N]��{T�5��|�?Ȥ�^V[^+a"��*B�l{���ح���{�x{ ;���=�B��T��c(-����Ӿ�~	�Im<��h�q	�
Z;�L=2�be͜X�PyS]��d��!߳o�	��B�29S��𥇩[9VZ�'ۛ�I��ԯ̬�'�#"�.�k]F�8v+>�1! =l�oW˴�;Æ�G��3Omv�]EC>P��kC�xKUǠ0��x�sNZk�*����+&>3U���E�K��6�+ˑ�����p�
a����Y/�uWk������d	wqaB���AO)1�*Ջ��}�1��Ȕ�x�66�`�� w>/�I�����y��T�"XR���^e�����gJ�p���U4}L�C���8�͝�q�]	�Ұ��ؘ(�?FX?��~hV�>8Ь�@�0��A������T]W�-0��K2�� ���pA	(�����כ�F����ן��lV@��-�\��N�:>PYI#_��[��sjo�.fj�i3�Ġ���ZHPGw?zt�d ���\S��:�:*彍��۫���i$l,J�%�a�_�)B�Qf!�o�KQ�m�~0Q ��Z��DS@������!�B6��2%���+��ª�\�T:sk`ux���l�Cm�8nW����q^�b���$@Z #9��1�Yۜ���^"�پ����1��R�&W@�j~��E�M���f��<z����ˁ��h����򍊑��sɓ����א�!�ֈ����������;d���rD�-�h�$��!�l__^3r��0��z(�ʇ��>4k[�9����E��d� <br{�������2�2�TIj�Wx���V.T�r�X]t���M��<������^odߞ�~쐃|�,=�^��A�Xn�{�+#+��S��#��q@u�#��� #��A+��� 1�O#Em�W�x���t\ĈUFL����X:FX�1��D�Jq�H�FuU2ti��%�V_H�]=z���+b.���n*ׅ���8�9��P�_��O@b&4��:�+̭4�&��c�U ��E q����N]9T�m��4�Qv��UC�j�դ�!kfY�Qx�;'18�0�)^��len4��>��&�]���s#���p(7�H]�r�1m�I��Ğ�z�3b�M9�(�Պ��A_����5"VWwـ�%s��x���ݹ�Z��-����F��"_.�#�NxpЈ�x[v�B!'�yp1Nl�>hJU��}윒R�K^�����D�s����q�c��qo��-+���T/_��m���֌Nc�B�����mBL��%c�AF� �������|��^
�U,r�����(\ m���!{ӏ������'O9X�����]�z���ݙg��{|����$�I�S��D�� �a�ནGK��'��-��3���8_yEp��3�/��q��Bg-�9KL,��>�O�T�l�+���g��l)g�$U�}��rL@�F~L%�M�{�b���=�C!jo�����Z���1�=;��I�1{%��;*�����钆"4E�\T�=s?6���t�>m3\�sG"2稛� ��~�3�<o�"�ڷH���ܸ�� ڊ�MG5���������������$
�+^�	M��k��Ȥ�3xKnߐ�@1�Ft���{.���W'��B�Vʧ].���Q��j�ԯ�8*��YAn��}m�AG�1I�����Wށ�a�^M>3%%pJ��2�;�B�ǰ4��JjS�b��eѩ��]K"F|6Tq�s���k{�xо���7��?YI�& ��/�'ܐ�2-��ۺ��[	�,{�mݛ�>�`���%��e^;��K��|��e����&33"V����~k��x}9�͵}�m�H*��lHP���ݦ��؍L;�Ħ��[���ޝ0�Z3��S�Dco	����Ġc��DG��u]��J�V��I<����jK�^uM��+(�G�E���K?2��qǸEFK��և	(pp�g�\�R��\�8�80v�]��[��HRp�~�E�������ڲ�C��q�3�GZ����)�秺�y�:C5��"'>8���EM��YM0 V%c���ʭ�����k�����DSE����j�"�va���w<�-��.�>�+���^�>�o�1�k^�����GjG��l��6� �6zQ}#�F�X��}����T�z������"_Dk�CK�v�q�6_����F�F\��s21o�d7�]xڔYP�#���1�՟1D���]Q9�U���c֌⡽8^��9��(����\/��s�����0���a9���Ps����r������U�ZA0��o�ോ�������|�	������q�v:鯸8*]�2��Q3����*=Bp;>Zb���͂NM|����MXn�6,�<�_JK6$��b�d��w'%8��Ob �?��\���}�d���8�A�=�,��T�l� �iۛ���7g�k�˭��o���"+qe�����Q���~y�SH%8��"�]�X���&'#m����B��_�+�\�G-9�0��>�$�9�3u6���k��|u93](�/���;�p<�@�eT]��]�*��?;�g�<-^��I;@�rwr@��M�(��X�[�E�F�SVT]�m�v��]/�$P���D��5J3]{9�5롋�ѾV3��*�J��{=�~�i�B���u�7r vt��_��n�H��O9V��̩�f�݆�Sۣ��ec[�A�!?W��LꋖӄP�z�Auz0/{�9JC�8"b�9�6>ի�3���w\bG��m\K�	�}P��?�t�f�;O�N�F����� x�v�ڥ5�`�Rz����+@K]gJ:����4��&��I�_ A.s�{6&�!&��-�Ȕ��d��i��#͛.�-���&�f�� ��_}a�3h����wE�,�3j�d;)S��|�&W:c�T5���1�̳Z{�š�ʛ��/�"���e��E־K�(��F���J7Jl �ʈKf�t	^��o�B������ �yt/�Z�C���R�Γ�h��نF�ˋ�6�`g>:w��i��o,*���N�*�*`ǰ�Q��` '_���������{���	#CN5�>=�N�ex�\�7j�}�AD�:}ѷ�+�2�%We�7Bqى�RW�]W*M�(φ\��oC��������=wƉc�X+�fbZ�z�b����ȓK���ס�N�Ԁ�uM�˘e�G���l̷?�U�mL�����y�Z�L���-�؏�BV%3�*�ѹ�a����u�0q�0ޟ�<�a���˄�/���@�#2/�8�X�^�p�0)�t���y�yq�`��9dF�R��3�ڟ���	��=�ʀ�AK���6�@�E�9����Aӱ/����l(��ᢙ�d�:�\`>	o�A�U�V$Ҕo���tj����g2���qT�h��:�z'��l�fFd -&�y
R\�8e�?�9
J�]�4����o��W��#r�>L�S������5��0D皼�S�	s�Bk	��Bw6�v`��B��c����s��%����}}��lzp)���b$a��5d�v����Rz��Dv���O�?�3u��Frf6�kFx�l0-�*�'���$���znӇ %�^�ɺ�[(C�o�����i�h��c�{��iזu>���?:�6�z�"g:�p.\���=F������ȉ��"������ƭ��}��;�<��"�)7@(բ�$����@*V��m74ᓅ{=���I��@�����3QC�*)�مU��G�_c%�����1~.�yJ���U�?�͑���wE��-��8-����yR�j.���.������5�UR{�SbG���l��fޜ��ߣo+~n]ٶ���l��qYP��w�;���o�W�x=r��*�%��J@�C�?�𧅶�caj���!֒#����i��-\e~q��Δ���MV-QP��;ϻ_4�Y�-V����A3Ci��Xi�0�E_���|����Y�U�
��@7$�AD��j;�lO$��=�%�?�M.��ɑX
RD����^z�32��J�77?2�8ެ��R�.��PC����֤(q)옘<_f���r����].l���Tg	��x��I)T�K�y�M& ��Q����VBi�x॒ޘ�N�k�/�Q釿�N�C����75������X��](�;���<�Vn�v�?�;�ٝzWәs��������'"Ld�;�Y,�l���ˉd��\�`% U�Br���;�4��`O��#��Yg5H��Zu�"2S�7v`�E��΂�A10`Mj����"uG2����j��{��%v[��j;�g }���?;H�=��0��j7�J��������?\~ɢ(5����r�ٓ��4��<�
V��Rɾ�=����NZ��.2��lh���]N�!�����C:H���$i21s��}4Z}|G�_ܲ�]����?Mg�i�N.��נ{n5@��A����ILu�!�+;8����3ˎ���#�'���A�N�.W�Ճgly��2Ơ;�u��|v�H G��ʥ���,X�1\���2��}��	�$Sx�v�͹ef�8}eզ$p�r- �嶷�����s9�^/�9�N*�����A���x
?�~�f�x�V`n3y����+���ǣ�ڮ/_���F����^�������k�ǩ���;U'�(�{{�D}����n��C���M,�:/J�V!�@�h�i��9OY?��;�����O��'��2�8i����'��+�����L���mU���+q�'Og�8��%v���Qe�8�pK�ᬛ=�m4�����|N	m���ԋB�Fb����*��f�X,������x���8ƙ��u��U�W���f'�JG�:�G�*���F��2u�F���a���芔̬��}\�MnƲ�
�Ik��ݶx��Q�[��d^�|b��;����I;z-���2�ti��sѱ��p����0��6���l��)�A��>:��ѳj�n�fC��6�~vzi��KH<��[of��R�j3j�h��Q�Xčn���L8�ǔ�BaX[��;ϐY
�]�s�BgF��r�<Lnf�p!3�<Q�z2�mJ%{?QJ�Q�k	U+�vs�C����Ǵg��%z��:����M߲�2#�`A�L����$횑/���ma�@?��ɑ����!ɪ�r+9�0jKOUEl��Ą�^|�5�؄
p�;��|�����)V�Pe����[����x���d��O��x��b��N�R���ﲈ���P'G�a���f����	5��V�����+^q�*���tu�� �ϻ/}�ۺ�D�����nNk��1�jp	��Ț$_��i��y�n���zl�D��_1�r�ܲYT��%�e(9K��^ed����x ?w��ӽ�t�^���	�u/6�C�DCܻ6��Xz�q��ڼ����,�đqs�=|$��҈�[��W���W�k�|��t8�+� �)q�E��g\iu3��e�����!���F����7�7?�O��DU�jW ��J?�M��>�
"zHlt'�Can�
_@�4�IA!W#�9�\to�,r�+N���m�����P���'����6U�(C�10��q����%$v�Z�k����?pIv�|�g肃�`�3�q`;�c9e QQ�9n��׍]�89�o�F&ȩ^7��a��,�Dј٠�jP������*s��k�-\:�F��Vz+] [�-k��!�9]��5�||g�=�������ug/��=��`���Dr���m�׳��r�L3A��Y�� NW���T��MP�����Y��K������@�c�j��h�����ч��ϱ�qhel�ոV�J����;�
�,2g���z?���R�m�����d���| �tj�Afr 4iz1й�b|�9��H9
Ci�9X�'�[��"Hrʁ�D)��[���'ֿ�{��EN�s�#�nmy���͐U��G�>����� X�s�)�����>�@�jYf�c��؃B׭��*5�LP{�j� s�	j-��j�Yf/�� J�Y����>�^����V�Qбi��_��C����[��8	 �V��0)��W4gG�|����v�Y5����.�K���4����075�x�yn����M=�{��G�
*�HIa�/Z-"� ���VОY�Ym�LS� ������Qc1:����b_�����N��i�	(�<��J`�Xs���l��+��lk͏;�,�T�u���T �W~�S)Ӵ n{�����y��W���m���A�nṕ&��
�����ʀ����Q��*
W%���5�TRD������(HHw1�PC)"��9��s��{?�?�E�<g��Z{?�9�Q���m�i�3-�/����p!����ᾲ�!��Mԫ��;fq��N�?�1�˙%/���z0�;���д]2}��ήH���8�۳�^[�xWAK����ٟ�:�d��'gC�IX�Oq]��@���P/���~��Cw��<��j@r?}���qI�U0JG�z7*�u�8��a��Q<�I�\�r�3��"��TIG���%`�^Z������f��G��'r�;����~�u�+�O�v��g<"no�P�QC�����P�KLDx��F�W��Z�-w��ɻc�����d8�����v-":���aj4��Z.���?�U:H{]�S���&޶(�����3.�\a3��>���N��$.��a/z6�t5�z�EN�XU��&aY3�tC/}�_�9�+����)F�uW��sU���𹃓�ZanE��	�Z]��y�0���� �=<"%�Zk�����Q���Q=.�h����,��Ŀ��?�:��g?��� 
�-���Z7�H[�C��>���<�2�D���d�
�#/�ӸS��u�W��ˤ�T�q�G��$Ao�z6G\md#B#�6�l&S�T�-Z��A��`V�WD��+�3���[�.�y�X�#�Hl�"��v����"�8�q�"z��jk?��~�.�f�f~P��-�*y8BY����m�E��(?�L�	%��y��%��d���s��]:���CkS �v��c!�����rn����gF��2E�J��5s�g2�!Wk��A8���뗿�'�^���=�8	\��.�|���F�S��u�֍\�����,�UfE���&�a����Y�X)�v����_$h��w�r��� �-�u��{��Е��ɱ!��~Gn]2)�pټ�]b�Йi���q>��Q���UN�	Ug�ɱ�3���nP����}�(r[��9����¶tBx�������H�P�� |�#��h�<9+P�l����(]���M��6<�&���r�R�8+��cĽ���<��q_�"B�@��KMOO�5�+����KX���ݜ����,xG����"xZ?�_�v�����P�1�L��'t�n���G
aM��(O���q��\�����z�6#��������f~�-q����'R�G�w���3�`��0!I��� �����5���~�)��y��ێ	�Z^#�E˸��%�_��k�x�B�̗��C>T�~�rogk6��������ݭ��ǅ��Z�yp��G"[�i��0)�(%�4��ZB�]I�;jz&]�5	���m*�l$���ź��{����і��0�����i��H��?����@Ka;���Z�$��<p�V�<�������>q2 �J��`2�.���N-d��ҥ�t���������.~��uQ6��G�Q~ 7O|���7ż�h�:0$_��]1�t�`��w��_	����Ec����g�3��[*Ą�fb�Ib��O���(�z�qe�B7��1���1���!��D 3�a�������/�Ϸ�O��a��r�N�/waYt2}�¬��(v�	� o�Ϳ�r�Hl~��dQ\\ njA�����2l�0z4�р�y��_P��c����(���,��Wի�c��kss`�2�����K�$y�!^�����|":E�n�>�b��g�>=1:x#ۥ �ـ���x�<IIY�Ŷ��-8�PԻ�ט��.
9��RN }�)ͩ&1��F���uօ��n�����1u�b��q迌~�����h=�u�i=��,���OȢ'�Ѳ�>+��=��Y�x�ey��I�7;Vz�l��t%=����Q���|L-F�%�:~�H,�[��%�K㤃��?=̀O����\�]'}�5�����nzL\m�Q���=�0��Q��-5w1X�b5Y��ʶgpi?C���
z?��I}�g��_�;{� ���w����Sa>�B K�s�oPW�=͊~��CL{g�m��~AC=�}/�f�����np���i�5-4}|Q��pG�g�d�jZs^��ۤS=?��أ�+�mԨ��):L9�~�>:W��_��	$�}�WP܍|`zu��s�%.Vc�Lt~���lH�K���[a��Za������l#�qOJ׏��cdl��6p�
��l6����V=���dE`kq�W�v+���F��ɗ)/��-��W:�ˢ>Ua]}�=��߈����. ����D�G�Z��P�Ѯ���dMv���[=M���3����@��g%���~��Z���{ַq)(Z��
h�#����|��R=�k�J��(���*��d&fR��}������a{�8�5���R�x}�%��˸)��=�×PT�<��?�F7�C���S^B�*ب31%��"�i����Ti��J�c�nw�:�1c�� ����~�	bt�7�M��,���z,�7셁��3c
 )���3�|�������֕S��XG���2���8�:�L' �Vވq���#��8c��ɋ^ױ*Y h#�@�K����c4/\L/`��~~�@*d]'h�V�������@��b�ź��iS�^�N��z��6�̄��I�K�l;�_湀*3[Wvc�b�:%��*Mu����gg�C�T��s�|ڨ�uN��1ʣkG.!�'����}b䌇�\�f��I��sZ�ɧ��U�{$�a�͕�R'����_��nڹ2��~���ie�;�7<� ��!�0��Ԏ�*S��-��!��8n@�>��R�	��gip�+�4���N� �o�3��c�=���{8y�h*���*������e߿�d� ��K@��KF�r2��qE�(���f��J�P��&������#t\Z�}��Q��[�jx	+�AYu}�m
��;�Jd4�S��Y�:�8���>|� 4L:�4�y&V��y7K�A�F���Y��_�q٫����-uI��uLr��=FJC��7�����P�u(��7A��j���Z����м��!V�m^Ȁ� �F�ٳݎ4���~V��Eb3��x+}ǎ�A�=��_�/L�(kӻhxX�p�'��F�1��3<'c*��7�|�1��*�+��;�l�˿�}Ҹ��H�7�Uă���h?�i��gû)ᕅ�\���Yz�ߛ��t�� 7��qp<��VK�]tk�G���A�x�K_nR[,;�y�a��!�� ;��uȭ�S�!��]��ǁN�ue ���9 �ЏM�_�w����~Z�U�F��E�R¼�$�|4]�l�)��hV��cѪ|��O�j��x���Wl��;�o� 3�M��~�:�}���^�����0չ��vs����=�̈́��0f}�*�<q5�[1�-�YFUd@٬���ˆlʌ�Μ���U�^��.ܼ�� ���yȳ����	�y���'�1�}\���V?9�p6wqi}����aw�+_1�j�J֧�n��UU!�����<�ɧ�v����FW@Lf�G<��Ak{9�!�^�� Z&����g�P����<�zk�(o�ӿ��3K���
�����Y�^��Ex�������
��q)Cݞ%_l��X h=,��	�h��5���7 s��!q�l��v�x 5+T\e��c)���J<*��E6���z��\he~�V�X�H7�$y(�����Ou}1�΅x(�*���ڜ�Ax9и�4�����5���O�
q�8�"%�m2�~��'�om�M�ߍv�_}ոg%��o�3U�m}?�Z Z�X��

o�w!��� ���Ei�@A@`�������_9����ˎ�&z��5��)W���G�8G
�r���_��᥁<�:�um�� 5������Φ�y	��)RB�~�����f���ӟ�\xs&^�����1�A߉^����"�N/K웰��2���Ԋ�O�5���y�tqyM�5�S[9�=�N��٭�tm���h���2NK�~�����8��ׯ��.9N�i�#ݥ5+VK�7:�ê�`p}iw:��i����8���B�K=�5����
��}�I`%�C�
��.+洈[u�zJufi 9����j���R�槰Ӷ�|����Kz6�e�"5��X�)��X�zm�1�F7��|V�A�R�NZ��g@�Hf@5`�l�3_E����3S�O�hٱ��}�[���=�4?�UU� �Nf<�mVU��|��������т��J��ZW����Hmb�A��y���)Ν8a<�4�5�Z�iH[ɦ7 @�K��	�����q��!&���w�r^]p�|8����������'��p v�c|������W��6x�_���_M�Y�TN��g��k��RX���$�{v;Тa�u�{pH�G\���U�m��a�ݴҤO�y�׾��s'�䔥B45�Ϛ���<I �J�� U�
��0��x}읏kzdh|`drfƷʶf����½� 3�Xx�
8l�>zY����t�����@��z�3N�A����Y�{nFt��@bFU` SR?�1d���;��Z�!8��p�?̐���5��,��j��7��k=�d�/~��� n�RA�����*�������>`r0�lTQN4��xb��p�� ��z��k/OJ�Q:�Q=>=�v���i8@�K�E7��ی�..a�R�)e[R��B(�1�����)�����bk�\��_����*�+��61t���1�e�%� ��x+C��`t�������y2Ӹ{�R{�'����.1�扰�����I��~$3���2��]��K��s�Bzo4���ח��w�P��|Hb����6v�Hd���#��0���f��|x��'ʫKirc��۷N��e5s ��m7�aI<�'���$�9I�9�ҺW糺�`O�քJ.��~�x6�w���g�����8_Z,��ޢ ��y@�!���v��(.��7�|0ٳ�����t3*@n(�Eg�)ݱ�j{�׷�Ք�śI�e ��h.[��?��A^{|Z2�c-��I#��[Req��t���EP�<����d�>�jF�
�^iz8�,�,Z���NΉ3��ss�D̥�ENW�W�ͽ�~x�!��ؘM���a��䓎uCQ���ğ�H�|�h�K9��ٵ*͖���� �*��ݘ��*��=9�mѯ��[YMD1�a��?����D�7u���ݞ�g	:��)ҳ�d]�˼������\�a(�ߐ���Eb��$:y���ɟ3��dӃ6� �@��?"B�iXu0!��Y��$��l��Ѐ.T�.z�ELK���E����B߶�8��4!�̄��ՐCn�Oݗ�	'�9���r9�wȽ�=��|ݎ�}������
���i����[����j�cyx��-�m��e�I�j������a�
/Wg4j���8��8K!2g`�.-D5-���ժ4�T��5�[�&)��@�>ݎ�ji��m�/t���5G:H=�����pog�7��϶p�&4�H��V_X����s�>�~���I$!��l�YS� 2u�`�����v5~�?}0:��j��d��]�W�u51�w�����쌄�"�b�y<�H�Rey�_�1Q��q�dɓ)�#�3yfx�6#"��r5+t��̱��f.|�o��7�a�O�GRނ���V7|��Y?�u�$����]�g6E)gD�k�̿�u��9Ȣ���ޥ�+^W�f��I6$d�XN�e�B�,��g_P�Ud�{�����w��g��x��j��t(,�Yh����o_���k��mg��.ГB����E���}zF��`��<p��-���I��2iG�����L8��Y�¨ƽ\Y���4���c��qn���p���F���u�_qG�厀Yz����L��8h��MV8JD��1��.���=����Y����>_�����p�Z��wN�'��^�tΧ]�BcH��52-�%	̰z���f�Ftʕ m�ĳGj&�1J��R��g�;-	��p~h臟�?}j� G;��E���=bae>x�\^'PX�@�c����l�ŷZ�gǇ�<��hZ��e�)E�V�<�ϑٯ/�J�|�P��*�����'��ߧ!z�ٳ���R���:��)�o[<��~}�VT���ı�0�0���OIO���'�R����6��V��E����9<Ulx<W�����~T�f�fP��{��X�����%`{Y��\m�X�0��MNw��`A�@#`�f^݊xм=�4�hXʆ�ݔ�S�Ef�������&��ieIK�%�u���K�{��������Op٬�t��:�RaJ��hN�����Y�A˳���~&s�UE��DGOm��E��71���A��R!�r�g?�<OU�*fg�Kʫ��^�1���5�v�V��Bx����l����c��^�P�?���`��o��:M_�0r�l9�*B�Qz���ķ�(P���8����j%�~V%�|��6���zh3��b�ga�I�;�rt.Y�Tw{��q�|C���(�$��Y� _X�A��;|��M��v�u}Tߜ�q!#!�Yd=%�l?���kT.�e�x�I˨�"2���=�]�B�S�N�K7j{~��R�Js��{��������:S��e��iDK�#c)�͞����*7����Q�6�#1�HINFx:,$�9�.���	�j`�gM΀S�YF���u�oxQ~1���[QqA꾜'��=�O��͍k�On k%JNu<���*WK��M��c���.��(�cM������0���^Q-GR�Rv핃}l� �J}�^d�U4�M��A�P�R}�P(�dF�e��.��C�Т�äXV�����Y�L-��Mx�s'��'!Q�t�]E�<{{��GxN�^��BN6Q4�\g��,���1��gg�lrP��=>�,	�<xP�RWǐ�Sq�%yg~������x�y�,*��iD��b8��<�,�(���H�nL�)���蹞��K�̅�BĽ����k&�/��8`Rh��N��gN��ͻR�u�\K=��:R�x��̼<�P��#�^&����>$ �HG`p���/}Y��r���#H]�$ [w!�Y�%#�������0�
 �);����C��1�#�ao�
�~��.2%���n]�\�2h>�Ax{��n��4TU����fL����=;��o[�^b)�VE�	a��������whʹb+��f3�	M�f��$LBu�,yRBL"@�I<7���/Y�/�=en#i�'竉�~D��877�]�M+͖��;�!H��q�:���[{_�U�!��q��!��iE86���?�ʮड़.ʔ��1������!6|��$;<gNV��x[D]�@�fy�I;�����W(�$}ヨ��ȿ5`��+J�r�����qJ��>����\���7��B���L%18�f�%�������l��ɭ ��e:�.�?k;�^_�a�d0�]�5Y>���i_�B�j��IGl�t���v���p�-��Kv�(�j�_ɷ�·!�|Z�/�+�^�HX�L�W+��c�&��Ck�LV�:�Ph�u���@���ډ��T��F�D	8��
���˳J�����>��o{FnǬ�ȩ��*�y���uʓ�*���������~
X��p_�Jڻ�nc3��df��[K�ҰV���G�*�2^��S���cu��b��4�q�����@&U�AwK9��S�<��l�v�7^k�>լ&�j���e��.y}���K�)̎�����z�K����B:t?R"W����T�S�Y��aqB6p�f�u� �E��ܓ`��%�d����������S�i5� %5K��t��{b��꾂�s
z�1�cG9�G�H���u�P:�ILd�^/��+}�&�w�⑴�����76Ny���_�G�D"
���{cA�����)JHe�ښE��E�Nn��4k�7v|(r�~i:
A����͝¸a�E>�U�z�O�)]��f���d�(3C��F�OAu�Hʀl�ա��1�0����!�ooh������VO��rs���d�ʢ���:(��&�'J/�gr�c������Q�*-����H���|<}%$���>��PQC1i�<����*k����[�{	����g�d��1�C��\�*����M���S6�P��b\^���9�>�~�c�̫�G�Ê}�1��W�2��OB���:D��S�=�zt"�$�{w����.7~�H#��O��x�_��kУ�S��ګ��ԓ�&���L� #88 �|��:߿����'�#tdƤ��tb##7���^�9F�ȩ�h��'?A�Á�Y�3� �� m��ϒC�`h��^J�+a,7.7�[�6=���
_�r�1�1��6�a��li>���~kb��͛j�TV�ʹ�i�nl������̥�H�(\�k `�1���/�2ۊ��?�ؕ��=ü�Y�*]I����X�V��<<��o:�=R��ɥ �w��qm:�ž7CD�Go���yS�`]"�Uޚ�}^����5F�R��y�-��}9�`�����M��#;p��\9\��zz\�6���p5/1Lȉ��gNDjB�C�G5E^95�䔁����q��TW��dC�32Gnf0Hʎ�?,"��.��c��44�%���SG��g�'��_;V��*�g�$�>��>��������(U?e"�T�'
M�ì�@�B7�u-�;dVR��?��&�m���>̴�=�yɒc�V�幋phy<�>�����g�+��Q~�K�f�2�l!Ʋ����bl�ni�Rv����>A�:EVh���n��h�[�܍*;�C��h����Ͼ/r����TP�{T^@���I��:`]\��?�P�
eT�G�U�~�����L��~�.��! �TК���w_�S�ʴ�J6%+{��=�Lc���"g��=	��; 2N�O6}�N9Y�I�e?�����AhFG0��9�]dd�ڜ�z��n	�*r�}Cc)����R#��_������KӸ>��4泆����*���PA$Yި��c�@l�YQ9{J����k� z��US�X]*���b�G���cS&�JΟE�Q7�����(��MB��!&TPM$�>U�ďT��R@Q1"��������'Y%Ś�46�0�-�=����� ���ݓ�g#o=���9X7���Nj۸�O�'�(�'����ě���9\�����o�x���j��b���������5��P`� ���Xz����y�k�&ʵ��)'�Ŭa��ù(ޔD��KN�nT�K햋7�U6FY������s��`D�l,��%1`�R'N����|a3��Z�.�v3WkBg�n�V���%2���]AW���]z���Z.���J�����T�zO��H�����m*��%Ge���@�c��<�,�b��P�a���}��q~� �7���-��MdvJ�/b/e��H ��M�?(Φ������Q����Y]�`��k��p���K{>��;��<+��n�E�pu����>"�$�~�r��p/��I�Y}n�R�B�s��j
W;u�z��X��|�/�����O[2��;U�H�p�����a�V͠ AV�S��}��ۓq㮺jI����+PT�:z&�RC`��qL>a����e�Dx�a/W>2~�_��	��ڳʯy��>c��V�O��H��;ߊ��� $C�bo6� $́�j]�Ǭo�[�Sep��|w����MC�LM�EYػJ'���2u�P�c��⧟I��YY�,ڙ�R�B����u��6U!�����w ���E�|�q�59�!95����L�jj���a�	��w�a�Q��D�W����،��H)9��5	�9[��c1���ъ�.��g -��D0Zs��3�Y�����#JŁN����gWD	A�m^�Ī
�o�Gl�w�=}g��b�ղ�ћ��>ɓTd�U�8�?z�c=�&;"v��������|��O  ��Ж��MFe���}��Ϲ5�T��xiR�cI�:b���cb��J�ԸT���'<����9TP�x��q)���D���o� E��(���*�v�/uw��0���t��p��P����Os�2� �k�
 �U�٪��'GR�(�X�:V��3��ʆ�/��i]��ɏEY�hx6���3���Җ��F٣S����ɏ�B����o��˧̤a����z8�8�;�|����� կ�C��cDB)��yr])� QXu�԰E��?j�$:$�6Vݧ�w�ж��������'��@��4��5h0��
<\s�,�"�=�<�%��{@r4���5�N������H�.�ǐIJ ���.�lһ%?�͵��|��f]��Ĩ�K��8[@�Kq�Yl�%�ɂ!8϶���g�:pF�
��
о�Zw���3�N&ԕ�Mt"�a�r�#�0�P+�ME@�}��Ia=�˚���4ݟ�~�u�A��YG�'=I���@%�+Q�h����,�O�&�B�,ε��#����t���)��������~|h�^J�4���.Bx�MR��!���i�o�<�%;�K���q��d��>�T���,�
�jX4���}|+����5OhAb�񈷥.�@���4�G�B�u�-�
[�ξ���e��c%Ph�����)�T����S��홺Ӕ�/������4���c[��}'���Z�f%�l���\����彵���C9�Ȓ��`�x�c����kc��x�v�/�,��k7Yq=yņ��}S�1��t��C��f��^�o��J+��=��}�g~���T+���?�C�S�a��t��r���&^ۇ��Q�4�u�_�w��f�>ʯ��	V��f3|rJ���d���3�R����a�{�e���9{�E�����ܑo[�@�,�="��걺[D��]�Kk�]�Yt���S��糇v?m��{k�[�A�%f����t����рZfa�iyZ{tX��x�(=y_7�^����y��r�� �V�d�Z�.GIAQ�6C�(勯U���^�g���h\�Ҝ��Pg_�l��4F��mɵ�b��%�����i��jy�aQF����AC� x�I�	�A��U�^>�+�W���P�G&64ꂠ��&���]�����&J��j' �Φ�lreg�!�Ks�Md�Z='�CPK �E�N<��:�٦�`���]�nfc�&ﺥ���|�{Ub�4Q�@���j�%/���v�~bk�A���/��]:�S ��e��4}�B�4,�xJ��û}a��k�����;��j�q���K�5�^�Gw7�ݻ�58��g�w�h4�n�(���-���<K�C;�ˋ.u%5��:E�[���Q��S��1��8썵(�V��7��rg��{uKC�����+f3w��Re�k@_�����oj���)vtZP���w�+@n~��E�5Au�E����]�s2:��|� �e����T�>`Є��t!��L��4o��WT Qrm�h�^V���<�6)�M!����j{ud�u0Kf��bW%���\r��� �@�=�|��M������YC;����G?:���VN����
�r��>}6���XNPY �4���˓����(J]THs�zN��{#�_��w���Um#d�X+��-� �:�v�$Iw��\a�0m��!�]���
���%_y����C	��a`kSF�m�/l�8:��!��9����2�I�������]"�?��"�)����"i�j�M����l���]7S�>�� �r��� �*�] ��_���coaܯ܊eiʟ�,1��Yn�c��3�����gL���R�%���,�z��r��0&� .��<Q�~��@k������y �Z�"o�n�C�yqHŏ���uT%@�n�T��v�G�'?�Ss������N�x�D ��� 7�*�Vg�X��jILt��z���׫F"��aJ�S �T*��yz9�WkC�Y���l�{!K��w6��nv�1��U�R��Z�]Uu�]�^X�I��[)��ݾh~�&�!��#@�so���ԕY��g�Ϻ�5R5�1��]E�l�������H��uH�t�5�=��R�rs^���p�h����T���61����i·K�B������n�Q��,�qҗL�dᰔ718��ۛ��n~�K�o�.`��>�QP�j���J	�6H���m��Gk��߆9ǰ����+i}x��i5+W�"gΧ�TL�	�
�gR5��/�K���/�"�5�(Q��'�������R1p���/�rL$3l[*2jv��$rF)5n����|~��|ﵶ4hx������޻���h�L�P��M+� J�����)1T&���5h�8���a�z�QQ��(rp��Ɵ���I�)Of��F�����ĿIU4g��.������<x�l�x>�s�����/Û�f%eo��}f�'/�E��V@������T9�K~2n��<�th�����H}����ܙ/y�b9e��c�H���s�����0Zꡚ�;N�|��^�L�mh�~�\�'`䢋/l{�ʻ�d�>��N�sPpK4*�3ˎ#��j����G���rɢ�lI�[�����N�đ4d�� :�ڢl��u&��r����� �
�X=�4�Wݜ*ѧ}Bhԭ�� �E��W��0��饡�r7i�k-_G����<����n}Z>��B�0��e�o���p��8��p�'3�J��I���V����+N?�;≭K��p�$�h/7�cs�dvp�N�U���Hb(+I�̙� KC��9����h�R���{8��3G�Ym|�.��,��H�Iz��Y��-�V˭!����꾃���k���#Hp0���P}iJu2����j���/��M���u~_ݖ�\�GLt���?�\ǕL��G(����>/?i�#�5#GRG	�.�Tw�<�螿���R�&]X���r|^T_��&{���hS���3@���f���c��O��R�崤I�)��;���F�'�|�SSB���
^p�Q�p��h���S_��D��;��!�;��s�2!�zߡ��l�;�t����ى���T�V6�p��#|�:Yo����m�>)_kB���k�\X�=!����*��,��ߡ^���	t�֢���kRuu�d 9�������R��w<��o�[j�F�c�����1�P�U릫��`n�<�t"ST��1��`Q���6�L~�R~y*�%����P���&���5�X:�Z�Vqkw��"�S�*�P�{K�!#0�����	���A8����;U泆k��s��)����%`���������oũ������q��ђ�s{rK�F7M�0I�n��vn�4�^���?�ׁl@tFe��+�Ŋ��T��*��>�%�+��n_mn��p��L��ס^u���g�~�-7^Lp�VD|��fM��£��2Ax]�n�e3≜ܲ^��������Rۡ�zzc��v	�;8�w$�&�zɹ�#}<m+H�l%�q����Q�I�����$I�8:pl���>b���ikq@y?�t�Ω�h�i��-�`Һn�d'
#tݩ��fc���HrM�=�1b�l�J��O׻49+�7ŭ��9_�q�&�C�o��+�*YK03�Np�bG.���&\��t+�y��7ۋ�"���PPP�p�����P�._�fc���tݲ�Z0�NK +�բ�����h�(�ԛ�Y�d)VF�hMY���1B�	N&#%mM���(%z^� �`��R+��x���ᄎ����Z��v2�C4�>qs��?�!�~#��ϳm�R�ڰ��/�Wl��V�����9L.p�=(!3�(1d5��6,�>��%�������L9.�o��Fp��s��RdG�$���R�A�d� ۠io����x�\�e�����$��`�ɑ�Z��q��vX$��/ܽ^S���HZ�r�M7{|�>�?$���g��z{��U�a����Ma�5J�yM#/{T�|X5vX�8s�l9׾��F����3���!������|�5��pz��2��˻���G��L���!@� �E���d]�j
F�i\˽Tx�@z?y"#�P'�V�Dr�A�"����ZZK��	��P�Oh�̡�6����s��{�r3��]�㧷��uG�Y��WK�\�C�p��6��)Gb���`w_��)��~`S�D�z�m�l��,�}.�Z?Xqpi�%>2L��6_� ��+KV,#K������o���7�˯Ҫ���n{!����H�ҜU}Bܐ���G�q��],>��F��e������n@��/'��Եg�~4�
������䊥�`�V�u7��
���QF|	?�Ûl���h�����/v�1���ox�6N�<Q��P�s#j�l�|�ܰ)˘�O"Vs�We�f ���Sf�շ�h�r�a�Ks@�3���2�X/#�ܞs==4j��y�4)qimq����	t�w���������p���n7�}��4����=�ᒊ�5	��4�RXZ���h�ެSh6��fʅ�C���;��[t~�Ī.�}���[�AB�JƓ�vG���=�P��F"avq�b��;�u���\"�Y��d���$�l�}sXK:��>Z �bT_b�:窇�F��p��H�?]�_ۋ�}�����G͞nJVX]�Q�/�Zfe�|Z��������+%�M��w�݅�}� B�C�Ն�}	�4=S��r]��C����$��������q��J{�Yb�������Tl�q��\�$V��u����\}5�+�K���uh��+��(U��B�R��Wj-��(�ä@�\FL. 8�vY~��������^����aA8kWH=���� ��t�y����W]?�0.�4]���1�U��Y��
1q���5�g� ����%�Ҹ��8�q�:�����*��^(,_-����p^b�P�e�/C��t���b&��V�kڢ��?��!��L777�iJiq�\���	DV����w�W3��� ﰑa��O,{�I���I�*@O0�~���I��#�7>����Tͨ�h��d��vi�����+���N�֍�%� _��ˠ�Q }S;D^��^)=y��!�%MY�[��Q�Y�)��=�cE�g-��+H\�{.�v�_��˓PZpZ���z����]{�1�����LI�-���]#�fYJ�t�����{[����VM�!@��|�mu�uf>�:Fɏ���ZoZ��+O<�B���E3w	>�1�v�	[	�����K�1����pz��wmyT�F�m�{;B�өׂ'�d-?������i��C�w�i��V�	��N�T�;�$H
J$��cP��3%ˬo�f�\�?]MqyA
���s��-�#��hC0�|KWy����(��#-�Y�� w���)��Q��P�����,��QP���	���YT�,�`���p��;=��?�J�EQu1�
2�E2��Z�2�ֹjR�W]Wm���A3�QZ!�\q/�a�>�HE�2uuX6g�Q���ִ�4r�]PՏ�G�p�qH��4��{?K�� ��T��TQ ����#\z4ׅp�<�Ѡ�����̠$�wV��cy�f�g[����"*I���(�(�>�aj|�gؠ*C���P�,u��_!�^��T�U�͟��?�+&&Z�䚳^9O~����<���`��5y�B_ -<���૨�E^�v�7-%����p��5�,��x�,m�?��	��;��G_b�����ʳ6����4���۽9�%��iCq�,Ν�x�G���$4�Uڸ]D]0ݢ�%z�e#FQR�-��nm��>5Q�rjq"�(�d�P3��ld^~�d#�1�:�9R�c�<.;vjjF��6�{�R�I��aɔE[��8'VBn�
��k�����a�U�#ul�����u��,߰e�M,�����UvO��"×tCk� ���¬��"�;��!K"���:�	c���W�Ĵ�-�:%�HW۽G�0)�����,'�-Rqx	h~
0���I%����k�{8�y]��e��r孲B��K����>/HYZ��DS
C �&�)z�N��l�Zih#�ޏ�U$� ^cmj���TN�'��w T�.y���d괹k<���SSĔ>��L�I�La�I%am4��ު��6�PA�f��K�u�>���pEG���Ϡ�{��H��KI ]�w��;Ǔ��~!���.�lo�3\O�Ͽ3�x*0�������K'�fH��D��	Y�r�S�f��� X�D��:n2W~����=�uBڮz�8x "�V�%G����+K�@�e�x���ͫI��7-H��'�]P0�,���@EkY����7�?��,��0�Qr�����2@7m���n�B����zVm�T)��dQ�M').�k\���;\'��n�[e�fa����,2<A�,uӦY��X!n(o�Pxw߽o#1�����A"P��u�InL\���.�6����ʜ���o?\؅E�
[K�a�'3�������v�289���Y#�����'fI�(C�<����T�#���rԜ"�8 k�����%n���{ޣ��{`�ϱ�]	n��˨c�:ol�2*g���y��}֨=h{֌�"�6w&���2��w>��H���$�k�����c?#��>�����}p���j���找v��-��)�y��-B�QZ��{�X�V�&_��� Y�Y�C��?âx(]mXFr���/{�.R��B)aH�b��rV]�����kT��3��D���[��MU�b��ŉ6�ʱ�|���٧6��׵�����lU��j�a��<<9H޹��ړ��[]��k�K/?�g�W?� �9��<��Rv��u�+k�o�Lx.�X>6��w�5�g9��a%�U2�4�s1�},dZ��:M����&J�E��zlӮbI����7�G�ֳ���7۶�@'ݯ��Ul�?;�ݓ�hl4�"�h~ʝ�4j�q�(Z�q��yXPN���&�!p�}�U���X��ٜ���[�)�/�ӿ���[�ve��������v~^r��C0"I�K�t>�9�����U���i�l�HJ�M�P�����I���dC��zT��@�8@:̭J}���X�c�"չ���o_:7�0"��h�qѶ�:�1f^w�R�i����(!�1:s�5�j��h�)�g��x�c�e��I���Ŏ����h�#Kp�G[ 4��c͡4v!�.:��
����ќ�r�aOs��R1����X�k����\F���v�W��Qr���Ob˷SN��Ngʈf��^��������C߶0a^u1 �6@�;�Y���βJ1�6���5�u���jKCc�	��2�M� ��|���X���(n�s0���0�gi��qE�������t~{z�X�N���U�{�k C�H���4o��Uu�mq�NP��f)p�OdXs�@����E��Η6�F��CK)��*Fџ������=���/ZB��DO��A����}"�{e�	���0D�����=��;3����߻�͚���֜����g?�{�3�[��8@�Ѹ��N�����\;󈈂,��n�}ZA�L}G����:� �~�/`���Wө6�h4�z��Y�K�p!��7�SE�����P����B�٦c0��R�]����D<����j�9O�J��a�蝥8>�iG�t���k��"Ü���ln����AC��M��kdG��L��+��������M'�i�Ñ܊*�OR��i�64���	�.�;q1|͖SV��gM
�ufKi�E)�����\�|ٗ��C��!���My�o��)-_%���w2��N�)r�Q����n�!�I�5v)��O��ۓ%���|췮�ܺ�4R�bm(]�%�ta1;���� �;�{~F�1�v���*���P���g'k���9jAK��jr��l�;�eN[�E�9��9&���x��T�[EiN����РG��b�Hs��-���1�Al�:���Or��L����V�o�l~fx�ὄ�e��UG�����������P��Y�7�������}n����p�����Y5h�?�u.&Ӓ�b,x��A��`��E\&��)ZO�y�_w
6�i�<�� �J,F�9U@Ǚ��A;q�x�j��u���L���3���C)Q�>����=ظ�vE0��ei5�VA2�9b�5a�b��L��
%��A'R&��}iM�h��z@�e��@��@�[�,��#KV;Dd�%+��Ľ�z����t� W�uuUi�y�C=Ck:����sj�vd:-�{4���t�7�p��S�2�R���szM�'0�~��h�j�$�U��&�hA,&��7�,;T /Eq�O�`��k[y���0%`�2�gf���[�_y������w�����v0�\+������ۺ���<̃֠���	Ʃ�U3���Pv�w�Qd�&�E�q���� �Z�� ��"b��L4��@t<��&,���# �ܡ�o�5X���Au�2�-�b�?��P�����¦�W��1�pxXb��ޣ��-�`�BteX�oZQ��Q�87;;G�i*�~���w�ab���b��}���C(`�ؼϕa;iO�O����s!�,J�`c����m�B���Y�� +��?�a�K�Q(Ts���(�����֪m�қ`3A�ȯN�Ϟt�̩Ҧ�&����P]:��X�w�2/ �`��?.d{oH����Q_�Ť���b��q��8m���b�a~�g�3�Je)�
�,��`&�@+�NB�%e}�bu>����_�]|�0-1��K������K#��$�!s�kk��؝���뎏H�/UVZSO�`+�u�n��h�;�-�^�}#6�Lg!_z��^QB��5*!���[&�:f�e�]�%�a�m��.E��C�����|��x��@�DJ�3Gh�}�^�GL�S���WJ��\�[)�<v���&���U���;8`u{մ���c
ω1��6��אs�l����˧B��
xTM���SQ����KS��	�PJay��>�ߟ���q��L4��U�E�\� ��.� ��jqJCy%�c���"mfj�~9��%^w��#�q#�a⹻�.! ���|>�T�U!��mI@Z��Q�|���IB�~o$Z����uQ�ޗ�Fו�MfqsY4���Р�c5�Dw���O*�	E?nb�k���[�{ٗ��7��{��tuU�՘'�ߢ9}��A=�=��Յ;�,"���N�z�@0���λR�u�$����5��h�1{.���Z#��5ź�j���V��z���d�d��++'�,��K9c`�?_��]n俌��Ւ�L�ƝƸ�gu���}c��r*q���f��k�e�u�@[� ��!��S��!՚�T�wT
|�*�;Wx&�.cb�1J�k�>y����f�N��~]ʤ�&�z��հ��P<��i K=�W��{v�{�_5g(9�&�6��a?�˗��|?�kɣ�v��jbQ=�L	��2���׽J�]6a���.��E�v��CP��-��J�v_>�ݢIh����1��0��Ԯ�K���EJ���T��(כg�'4��۝��_���m�"�V��мʆ=f��+��e�ຼ�R���F��"5�K��2�2r}�͸�G��y��E1�S9��˘�T���jR��z�e4�2;G�N]�3'99'���?��gSf����� '���h6�{��t�ϺD�	RIO�i@���CS%.|�M����bL�s|�w����!����s�K�h�I��l��K�}E��H71V>̕��u������E~�(2� 'ac���j�(>�H5���1���OJ�����+�º_^�1��%9���@%;}A>�-7�@ �Z��?3�p�SI��.�n��:Ԕ��*u��H���+O._�<Qo�&�i�����K���>-D��Nr�`�'�V��>ޑ�#��7˖��b���s�ð�����<z%��CΙu'��,yV�b!x,e��+���Vo,�ǳ~Y,K���@��*}�g�( �ȷ*�:�\_��5�>����٦�p��;�[��U<�n3cתE�C��
�ēr%Hn[ոN�/�|�s����E����H��C�USM�lI§%z:_gQB��|B���b)��p������X�[{���3�3Q�U҄���o}�%X�I�L�^�@�l���w�a"#����sU^3����a`;R0!��ٶ�2��+%�5B6�w¬N�4�;<҇���þ�s��-T�+��t����,�%N)�E�O���<�
�ؒd���6�̽��ᶽ��rn�!��:]���W�}�p��6j	5��&��� Bs_�����̃�ً�����|����&쎏�ܼV|z=�>�n^�@:s���mx"���=��U�F�������*�^�,�d��Tȧ�p6sHC�ښ�J�j��c��P��_H7n��Mo�ؐ��m��<�N0�-���()����o�[4HI��Ǌ��L��=Wj�[<|�����	��K� 
�ֽg���æ�tE�R��|������\�o�7�7���}�läRP�0Ffa`*��aǷ<'�H�$��D���}^��@T��Ka�{��t�kBK9���+���`j��JRtm*�<�y��Z��d��uJP0�f�ペ�Ⴍ��L�o)�b��Ht�w3���#x]������dj��԰7lP�&�۞�^�Uu5��}�Q��gi����C��,�V����~�`���xv��;%(q�����Z*���'��:�Mps:wz���	ww��3�kXb��櫎21bJ�w��]&�"��I��VYx�/Kè:v�߾/w��V]��(����뉣o߸\)���*��=�Fɟ�L���.Mؤ���N�Y*����\0��l��P�a�Ob=A��چA��A�<�?ͻ���fU�5_0˷�Ȭ\d��m;(w��|ifc��R3���a�4���4I�K.�Ʌ��݄O�%���q�~� �v�~��ܟL��|�ǜx_����y���L�m��_
By��btN�=¯���� d*��V\5m�n��mS9,)�%�y�alXm2��G0�A�A��b�<ޝ�(��3�/~��� ���J���/`�������uO�T�%*:�E��f��bGEOD����*�B"��7��r�J���\�7P����t�Yk8\W=��ܾ�+����l�r��m�*��ꚟg&>�9�����%&5Iw���RV��b��3z&9X^&t{m2�K$��o���m���ec����r����cD D�����C/���5H��*W4�,!�S�!�Y8yP]}��QV��!�U���%$�w�R���0��-9�$8���)ǰ�����f�ꍹ$�H�����a+��zҫ�s_3J�?�B��==��QJno@K���3��q��̃A��GG�V�j_��;���I�F	l�r�G�М�3���I�Xw ^G��yQvqE�M ��>��T�G���ݕ~;�����Z�Z�^�����'�J��1S�k���Q�Yu�|_иp��d7' H�WT�ڹ��﫪�F��5�d�������6¢��ӵ����<p�\W��|&�5�T*N�v[�b�V\_���O��h�l�O8ܶ- �%t,Zt	�[X+���v�����\?�= �u�(�T������S�4-��~�+^ա��~�����ctO�ſ��lc�z���JJ�L��kEO.v�����#<���u��$���ݚ����O��G�ie_���?�5�|�*��.�{d�[�O0��b���;5H�WH�	1��w�]�'�l�ȷW���kI�0���'�>2Qd�y�����ǒY��y���rD*��<~v�� ����Cd�#ث�f&rb�Y0?�hL�ި�����<f�����?,%n�����ߵ&��-�iAz-M"1%�x��8DV� �m�nJ�F�á����o������N8��f�]�Mk7_R/z��Z{��͕Fx�������b&r��+��U��ǽ�z�ܥ-�'u܉��Vs	˿�MƬ�&�pYl%G1���cJ���L��	����l����W�sR���D������N9J��㬹� ���)��z��=n	r�t6�&|�=�.��n� �ͬw���Z��*�uz�j�"qK�v���M�h��@X�ǽ�׵�o�TV�szZ]R)W�8��,��TWy<��;e8Uz��W':��!�P��0�hgۇ�*R�EI��F�/n��̖Z����K�N0���ğ}�ma��R��at5~$y�7��s��Eq���4��_����.OE�<��8E��YJ�nȣ\�D57�k�W|�h����P��=�J��PV���:Keh�T��6�TS�7 �����/���פ��*��rfPi�L��l��{�^\�	c�2mour�Ѱ���M]I�3B�ϋ&�!?��h#�&!c��e*��OgD�4^�J�����������$�jW��$p�љ�%���ü3�n-��]�mq�IRLUQ�N�<8q�#�̈́���_��_���<~��M
��l��_�C(���7�>�V�0��*?�׷g%re���6������ߍ��3�"��B� }�Hb�����a��Ǒ��z�������EY���&��`��ٖ���}̊:-�LƫyH�`��{C�l�_�׽��e�8�G(�0jSsBto���jk�	D!��=���]��7X���z��9���f?�fw�ɯ�-��B��tƐ���v�ߨ�;��ڪ��IB-�*�I"��AJ�&�r��6������oJ�ZL#�[~�C�/�̕{r{�<�/�|U*���\��'��������j=�@_�����0����ܰ�e.BC
?����H��4i��M��S��X�f�82���̺�6q���>]�v�$�-����X�]�U^�����|��d�z�I�|�}�Uw�����W&	�X�%�w���#6QlˊK�t�[Kƻr�����u��Ԉ�m��F��kZ��t ��E�ʐ_�A�a�AA�7���Ӹ4����~ޑF����a������#7��aߔ�x��z������(�-�tl�7���`���,�b��P���F1慭�b,5�ݳ�>��O�7FڏWV�S���\ZXX�0�#��"*��~��ƙ|��x+���,\Æ�c�K�Z��&׸�jX�]����� �_MԟM2�_��#�u��Xث�ǆK,
�����wO�HmH|���Jw��rf�����oe�}��Ȭ(���xJ�hM�����$J"��aч8�<\�Sؽ��.�9nl1X���@df��o&.���l���{��Pq�6�2����Gx
���n��&�����1(J�0���1Qlu���l:�e(��ak)*���&Q���#_ӁEǂV�?�\��Э��
��9Y�~=�p�l���q^]��~�az������dvT?��,x/!���/��<��1UUcee�v^$*�[��X����j]Xۉ#~-%תJ��I79�պ��Z=�.!�w���K3�Xy���y� ���/��un�Y\���&���X�Y�4E�����cu8�-{�`S9�������Z6S9�����3��S.U}���݉y�	z�^��k�`)��8�
>�ޚ�?��m��~��������@A�k�<�U�5+�1�*�=#D�}���!�,�8�s|�i�D��VC��j�ԞUt����݌����`�^��s�� YOY`;K�pФ�CN&@sAt�%@�5� �;~��DZ�iI;�����Ӻe���g��{�N�S�[^��x�d.��LDkY���M�\��>�������qN���&8>X����V���T@$�٪Ȃ��O�7KJK��Y������
����������1��\�����h���Fգ�v�[S|�J���j�U�����Enf�G@i�d��ԃ�ݽ(��J�^pF9>�L�>�2�eJ�=�<���ka�]�J;l�dK�R�\�Yb!�a� ?Ĺ/__����UӜ<y''ϣ��(v��j�є����^�O� � �)�ég̚��g��Q)_/�m��y�]u�mT�A�ˡ�	bQ�����u{yޞN�|�mS�d���꾋SP|H�0AJ6<̴��Q4'gpP���nj��mL���I�`�=Ɛ�ͣŖvR��"��`Z�n�M�v��od\�fS��0>��<�I'<�����I��� ����#��<(�~=����w[Z蒰���ܳ�a_��9��]ɞ���wr���b���^J�,���l}��z��:1�i+��t9��qdq�5L5��/*rk�ЗdhV���(�d�@�H4XLV��lQZgs
bE����>�}�=�����-��ѿ�F��6 ]�'����?���Nv���~W�tz��֛�}ˋ����'Y6���o�Ȁ�fS����?����s����8��r�غBi���q�B@��@���\�;�n,Ɏr\���W��K7}����,�~���Z˛\m%����g��,�Cwsu����^Y�����9�8pc�N}��żN�-[�r�����L�BE�;y���"�
PX���B$������Q.��6�6��+�zi��.�+˙3�g�+��Y{F�/0�� �Z��"GLt�����_����ln�O�Ξy֯+O%���}��[�>%AQ�����ٱ2��L���MI
pYC�sȻ���Δ�S�m�[O� ;j�bD}����6-_|����`�Jû�ire�
�X�z�eQN�`��c/���=X�)�9��Z#�֤A�����o
���zs+�e���D;�0�t.������'3�49K���+t�Ţt`%�Q���ZO~P �f��k��R
u�u�M�W�i./f��4�+�"5CY>��DۉM�B����4g��G����m &�QVX5$~�~|�ָ�X�y�N�)�L�ԂF���̨��n8g�o��U����1�҆l���<���E�m^8O�^��m�i}#n�ڛ���Z1ڬ�9��:�4B�b�r8�֐�7�ˡGv�sT�-(�U���(l���\�
�'I�UɬoO*��ҭ��q��gU��M�b]v�Ӟ[p~�b�@�r� �C�QK�j��X�4q�Dj�R��6�*%2�$H-�/��*�F�����+d�_�fS���dy`%����O�wY�X�ų��9N]�UYI'.�zeE�����ӱWڅ���p6�G ��L@���w�]Y��o�r�(\?f�.t�eq�2�]'K��[������s��%�_~�Q��<�R��nU+�74!�em��Cp�ⅰw���j)}��/ňy���TI�>	��]y��?�(�E�$�pK��ؑ\n�I����[bEyW4��,�z{
'b�Z�╔��z�;5�JԙMN��6�J �ejV>o��&���#]@q���r��6�I���_J��H�{���b���PӍ��W��*�Ӯ	1�4mVz�e��ë�o� i2m��,ߡY���x s�kD���]︪�`���W���*�^�-��0�F�N�CV���_E�!~�m�U.�3��^exU�nA䟸a�C��Qt$em�}�c�V���N�SG�Keeb�K��n��ʩd��핗y�,�O+G:^�G��$Q��s����Nǉ�U�)���(��#1���*��H s5!�=}�{C� Z�Z�R�<d6� m�J h�A���՗�T���:nؿ!L�w��>�-2����d�.î'+���A;M�o�C�'��*�|��m:����a��S��,���IC�����xNR̔]R�n��aE�� +��|�!!u\�wv���2���b����Yv:��/���u/�#v���;S�T���̇�<[�?/[Z�v��@	�����k.�m
�N[j>�d!F�P���`�aܠ���W1^�H�>&�{5�1C�p);E������g Y�\&�r~F���x�}�Kc]ڢ~J�N�X<���Qs��g{�/����TGg����}ӡ7~؟�a����F���M���DK�:W}�v��kpM[�w[�Y��B�&�7����V��)#{�\�����%Lg�$��d����	)gZ��+O.���N�� �訽��\>5�Z>��RG�RYpN�@����mv���k��Hbc��Δ$����(��7�X�P$�����fzs��U���z��CW�ݵ�f�Q��~ܦLE�TV������oUcl'ΧnWk:��$�eq�����5���ɴ��T��:�䊺�s���3ފk&�F"~�{�{����V��>|���1j)��7fP\=���Y]!������y>����~���I����b��=:�s���9�2���A:�ؓ��W�l��wܭ�]�S�i��}��.՞��Q�+������3j�&��Q�N�_E�̟)ڄ��ǫ�{����m�.ͭ���D�]���DE0��"�N�I���L�Y�<b��!��¯�S��y0���'��L��ލ���^�Ma}���5'�j��M�����kw��~����I�M���qg?a���Q��4��|'Lzwn�`�{��|��<;ۀ؉y��C���(��w����YxL�Z|Ǫ������òjֆ�"�ۯ�ϖ;��P��C<s�����uu&ԕ|�6�πƲ��q��P�����y��P��w�e7���`5Jes^�;���m2�T��j;;������b^����I�^�ގ������H,��/z��,3��I�%$?�+K(�~���{3=	@P��ю�� �w[�_��o �s�u>��DM���U��<3j�!t�g���d��29���YG޾�/�=����ek�6h/!����RpNN%��������5N�]m#H1��:�sD!&N��.��pc�?��^R��äH�S�!u��ABϦF芠w�����ɝ�L�o9�}e��9��iP~�x����7��wx�9�9@4��]��5�\Oh�'A*P"����h�c��)q�aH�y钲�Wl����})�[=��zMq��VJ*m�Ϲ�]t|PZUf���.�?ҥ�wb?�&����e���9/~~�faHLAge?�S�
hKZ����^9�":�)e��D@�vr�d�g��Q<L���p�>%����ø��v."��=��A�",̍0��uM¡i�UC�cɔ�~�ܤ������a�֏���W'�൷(c	�G7H2�B����S��Ki&l�}iwD=;栟Q��1���`8]5u�ޤYd1(\�T?�F�ȓRЈv�r�tS����O���1�X�1[y�5������}����5)���+;���Zk1n��)tN"�l�v����m�̧aʵ�[9r������;�ߞqr-��R6{G+Zq��ɢ�$�����\<֟��P��PK��:�kC���&}O�E ��=�[yQc�h��ǆ�]������C�n�O0��qR�����8们�3��Q��j�d�M�Rd𾦲���%>�0��E���]��y�<X�oc���n� >�9𥘱>Q��%���f�����`�O���������b	UJb��jd�VI�4)@�?���0xMo�ۙ%�~��x�
�0�ݲ��-_�\�<������y��J-��AQ5V6�Fs��-�d�U�e! ��x_��U�+"!y�t����$:J����K*���O�u�f�edul�%���o�z���C~C�L�~E"S�����cz�����	�E�/���	z�9_��c,rm-�	��lԘd�	|I��2�IĭǹNb�/.-)�H�ke�����!��b2���`��0{���`y�
�����NDx��s�-��XVƧϷ\8N��p���cNX����L�}sE�I���WlN�8�z�\`�����?��
G���G�ޝ'g�^����.g����|d�z8����}�V���<Y|�����<c���X��bo�$���hT�\���2��M��	y�^��V���O�w���Y",n��ts�U�A�n���m���dF�
��ۥ�.��	�mz��2��/��m,R��_<�m��K��9T�I�ٜ:�������S�-qR��������L�����3(0����P����;mN���U��G��j�o�bz�	�P_I���/�<�}���� X�E�o���楕ɝ�l�23��,f�~�'��<^����:r��G�]�u�2�k�6 �?̬WOl��K1�ђan�[c!�0,�� �J��	�c���T�B_l�]b:PZ��Aa�,;(���7��6��I�7��;<2��`:�:��#�$*����柝�0���ݮ���1��2��B���}&�m������GX�@' �V���gYMر�Vg������=mTe-�8Y�@$��w�w� ���W��I�\[]�=n[��y5)�K����5TrӘLXmWCU(�z���{~���b����?��n{F��b�/u�K��M?�T�7��ݓ3��<#TP]Qj� C����	��m�vCj\�©�F��{&���I�Fq�|��N���Ft�+�̙F����*+̦�i�Dt ��βNg	��u�N`V�_,>S��Q�:ߨ��)�SN���j�Kkf����%���زm���,��|�α\�@���`'���DJESr/��㬸�"e�|�'�����],�[*V!����ͦ�9���Kg��Su�3��F�3�!�-A�bG������O �4�o��� pPw��
�<J� ~|�ۑ�¦$���^���c��FX���T�Dd�U�����)M�"z��C�-��J��:&�0�F�������z�����<���Z��(>W�f�����$
6g2�y��4D���W�q߸�'�Z?t%Օ�"��� �s���2#(��&~B��ͻ�t�Xz�6�8u�����7G��OT���!�.�O��;��G��_0h��-�5��=�n��<�ӦB^��R�Xq�X#�C������@��@;�w5p�K��\p:���ixzy%K��~���=k�6�%�6�ib�~��T�����X��˗�ﾸ�򞎺`��~!Л���Et0n$��AL�G6��IƊ!f�G��?w#��Y>M�?�cӝ?\���ʩ+�M�,@���Y��J�{�m��1�C"e�r\��Og(��96�к�Jo�lŤD�9�H� ׆)7V��w]s�Rr#��n۩꟯�'��8��H�]�Z;
-���ҏ��a�r������������;����GYb�&gG$O��G#�g���$ ��ba����n��cO�/�k�<�mX�	yq�=��T��ә�}��������c�F2�K����bcm-�u�eA-���xD�p�|�-<}w�FU�a"@���4(�^��q*N[u�$�����J$F٥X��=����M�:8x>ZQE����Ǩ),lc�?u�����H拰�N*�a�t�s�t�c]/�2�t�}���88!�����O�	�c��TNn?E�<�`h�4�Yv��m^���h^�iL���a�XlH*���Ӿ�_�������蒝���u��+�j���Ot��O�C�Uc����`mG��w���'N���}�Α�|�R�t�N�Tj7"�7�m�+o5H^`�~H#,B��-���>��7��-1����6=��}Qg�J���]#�s��;�ִ��L�H���SQ'G�V�U� ��>�6����p�l	����X<�B8��7�H�8��h���
4�f�3�m���j��fڔY�c���6�V�e�'ǯ@N��W�7L�cA�O� S���`�)>�)��u��$��Q���C��|7�#�Ϭ�E d������nX�h���q��v���B�3��E�O��u�ylݧ�������S|��e,TZ�zPN,��lw{n˷��Pf&rf���nS��\+��--`���O �=ʎ��6r�0��B^���bb$��7|z���-�3�5��"��H���[ۗ���l���KQ�b��g���<{��y�Q��w^aUA^�׀���u@=e.s��>�o�q|Jr'��re�����B	�^#v��q����Db�K;�J�G�CLI_Xh����b1  hFw���%�dBb�\+��o���f�jQbn>�ޛ�����t@
�����.�g�;{N+�B�݄�lh$�?\��Q��VuAq���N�x[d>�ز�v�%up��������ˤ�.ͅ���ls]�4�mƛ?/��k%�E��T��f��yK� �?������0n\�n��r��!��(���yR����7�Ĉg~���a2����s�5먑�j�̧$-�?�]i��/���eQ�30�.����f�����麼�d�g"�ϲ����M�~{Wb
=t>P|��5� �̎7�ۯ�n0�m��;�+�[& �y`?�:ۻ@S�J��M@�gx{,�9چ�u��k�om��	�)��C ��e��Ϩ�,��҇���#.3��@,U��|@oNf[�TR��f��P>���~.��< lΞQ|�놋�M�,TvJ�Q���H���`�V����mg��"|i�ǃ�4��� }���x�`�gKZ3���f}��?�,s�㵋~��G��u�{d�no�&�wL.q��Rxp��@�%����t����t��2��ϓ#'��4�M.xŴ:�Z�]������]5��x�*���'do���v=��
��q�q�5(��m\/'�&;LB�HM��T`���󜏇w !<J�%���_�/�m���e�l�m�W��6_�x1I	��[�ls��F�e��*��0���?�8��wM� ��5CO~�4�_����P���:�J�����5�0�h-n��W&�>v#CȒFRT���FJV��:Τ 3Z�}�~�7�3�ܡcu���	G��&F��<7��jþ�d��	���!@�:�)İ�r�_��~�ָ��_�r�uw �F�u#ٜ,�(n��|�7I�xv�ʼoe�7���/��w�7{?�� se�9��0Sg6���`�pA�(������G��r���`�M."�g~�w��?�j�H���4�ۼm�J���L2F�"U!��]I�Q��5qj>/�$��9b�!���t|��,����@�Kj*H�4�j�\(����ܖ,q̠:?iN��V����e5��xh�������ve�N��S��߯6��f"�=(S���ӓL��z���3��<<Z��{�s�O5�7k����Y��J��[K�� �oJFL~涹rZ)�a�BL�ۖ/ct��)p֓p+gh�Iw`��+t�<�j�q��A��^���+�|J�;ĹO��M���%�VS��\;W0#:M���}�BF�Á0�
c����;6Co4M�� m/��F�#����:��<�5��KXl8�fb�Tj�4q��m�!�f8M���G��mJ��c|�'_H`�_�/'�OtAΦ6���}燥�����_}{����N.��.h>*�kI§eup���<��+�,�b�.�&~�z���o�>[%nu0���q&ƺ�GQ\^�l���k��N꿋`����,8�cOL>5���������������=��~R�.�Sѕ!��Q�Z��w�r�͟�T��K A%Di�v�ȸ����P�4O�e�)�Um�������A7e7���Z��Q�x���w�4������ן�L�cS��67��/�
o&��=�P��X�'*}���Ϩ���n�ʔЇ�	�v[�q����
cw�{1V"�Z'����=��U+��v*s�Eu,��`u��D��>��-����-<OQA�R���>�w���n$:�k[[��D����{�|
����ǅ^���`~��u�GU���(=�M�d�"����J�o�(e�v��y�6�G
�N�Iz��;�v=��~j��������et)1�,eI�<B�*ԁx`�3
F��PQ��#p�"b��_��Q��Bל���|i_�'d�E����:%��'|2�f�{�u��ӎ�t�1��J����s�5�����l��"�)C�K�5��'˪���M�s��to�D,���s��r?�!&���M��ڕ�_�>5�=�G�.���	�\��'�%L��o�`R���F�q��r�%�QI��7Jk�D���&�w���B���I��i�Jt�>P �mA���f]��^W���o=S��Sǧ3S������J�e��}�ނ�_���; (�M`M���?��?�,:p#j�Ika��Uu�{�� �`�G�xa��b���E*fJ� ��1>kZL�i8��Dr�5�2���;�6��&q'&��u���[�Y�;}�I~�GT�By=%1�����q���wO
]v�e����t8��x�H�^��F/�=9�&��~.|��͆�4�x����Q��4�p*y���(5�6S+Rx9�Yg��*fKp�m�=�����`�jquK�1P����şg����sE�)@'�h,���I_h��p��{3��	��{�"��n���6d�&r�k٭v=��X>D=V^b`��?�ƿ����(�"�ֺO���~��� �,�N2?O+�˓J�bL5$�r�|�}�#����=X_~S��̜ Mb�P�q]���]s�]�u7��������.�S����UP'
;�h"�M&{��}��Q�R�Ƀ�:l�� 
{^gC\-�n�}�F��Ӂ'3S�A�v�D�k���Ɨ�Nf�O�z=�1S-�X]��g���ӝB�`m6�6�C��S�}��E����NĵNoԢ.�z}M[�0�v�ݤ6�`sp�T�I��o#�yWB�&>rw���V51�2?t#���,�Q�Y'[C�x\Bn��+=֢�H �����~�}CD�ݛB�h�'��Q�1������_��v��Ф�������s37� ,r�^H�r)m����������Ӛ?������>�K���s�nr�޷䣈W�xő��v;���	�h)8�rX��Z��?9��y��U�OX��b��0�F�lF&��	n��X�	W��jt�t�`$#�G߆�	�]����=/�h��ʲ��]��fI[>@Pz?�:!�bF��ڍT\c����
7bm�$2��;��|�/������ș8a�U��U��*)�/���G�B�,uQ�s�H���5T>�5U d��!��Fv��/�0-�"P�{����$� ��6��]B&�u'+��)�����q�X|�Zxo�Ԋj
D��m��L(�`�.V@����5g�_���^�D؟��m���%��g3֛D�H#dWx~h��6ݼf�.\��v�W�c�-��,~�EU�>�WWC��0N0Co�sx��l���f�l}rI\b�0�l�,�&�AW�'�/`՛� {�*o�i 9��8j�����_�a��lJ+U���K&:���VA���<�S�lҴgB��Ƨ���l���K��k���N~y��D��5 W����6I}�@i�y�x�xŠ_ �L��x�^�U��˨?��HB�+zs{��̓�@�����~Y���c.2��Y���UllY��s���զS�<��=��xt�"c3����i��^Ƌ�l.�'�@T�p�������-|gެ1ߵ�"'��)n��V9�k�E�@d~��Z%4�=��_��2[��?"?1���Xy�1#����~j);�nV�6���ߎ&�H� ��r$��X?�����'�qҚ���v1����e��Ԙ�_��N�Ժ²�����[�@��~��~�s����%/���0\4m���C��khb�*x5�pR��	�י;�]wp_4h���(��VZ�-��������3G���-�'�`�*�(/W�:�J7�2�\�������[�<ֽ0w^�E�`j����랬��t��G��������d��p�yy�aS1h�_b|�ox��;t5�PE�n>��Sx{p�j ������V����f�5���ss���'��i��`��py�B��41�	oX;%�A������֥��I3�I��pv����,w;y{���0L��ؕS����'�w��zWCan�z�B����+�n���Ƒ����6K��=�o�u�Ko�=��k}�����1xq�R?+�E�<��6;���M�������}A���EGe����Ȳ����#������w��m� !A���&���0����z������R���b'�ͺr,m�8-s�������b��&��6��m��#��iA՛!>�D��mL�9�3��h"�Z��.E����n�����Ƀ�����e��^m̀h�0C����yB�G������h��q�v��q��ĩa6ԥ"u	�8-�A�rv��x�X�+ewE��W�����^�������<|'k�����%u��λ&i寂T�
{���Z���ƭӉ�23�\���jK����P����"�c�dR/=�ߜ�6T�6����$�%���ɔ���*���Aa��pY�!�!��)�K�ϟo=-bwf|�t��n�᭦�α���<��k�ʱ�c�x,��-��1'�����Ԍٴhu��G|�����ՙ>�>�A���h��FG�[���IsC���7��S�飭�ed�e��=!:?��躛�)����C�w�5u�m�Z�V�R"�
��"#�
����
**� �VA@��T�2e�A�=��V�����|���}��O��Gr�{\�u_�sN�3N_�M�'�[����Gܶ�ͤ��b �M�����Q���Ƀ�C��ov!��g�yt}�Q�sxo�oQ��;�˰���G�������8��uKFS;S[}����(ë�fPh���D��/��e��g^5�5.J3K�~�AP��P3�1��Q���gY2UVkZ�5N�G=8�>��]TXK|<��g}
�B}z$��R��{T)
|��7��\��o��k��-�c�7���P
j���[��vd.����~��֤��?����H1����2���8���]�kc&dwg����O8�?�:�(��/����T���v����7�����?Ӕn�nu�3<z7�SK�O'ӗ�"��&3���l�/�j���ƺO�k�@���'(��\U�
4W#	T���Mx�g�|zj��4uR�im���=�/�O�Ĩ+�}WMb,=n������*f&y=ƒ�]�."��o�ٽ��"�"٣����e�ј>�UU��'��o�k>0[�,8>�Rx�z�z�� �3v9�>:yu��|�.�]0yw��Mn�\�����X�7@}Oؖ��ʢ�?l��ڷ���e~���+4
�|ha>�Ac}�f�"��A����+`�_�:l�H'�'*�?K�GW����ڨq�"T��ff�F�*�.$.���a���?+nL5�p�OɌ��U�"�V!q�_O�����g����?��
v�����a��p���� 7��V�s�
�{������XI<�_�Q��-�)0���*Q��W�{��7�N�H��QP����(\�N.p�2���9����i�WiX@�6n�U��t:�BN�N��}�a��ċ�z��=�6�`��Z����|���&���k��`��ƞ��N�<N	��1�د�~��B9lDN�q�W��%�嬠A�e��qD�~��ÖW����[���F�\
���k���D���5������11�Ig������|�4J=�!*� h�IU�c���Q��4�B�`9���,��*�"�=�C�5,=c~[#���r�Av�r�t��-CPJ�n�!cqjG���o6�dV�D%���'���e���G�9����ŵ�	d>��~�0�u��k�M�Ŧ]]Z1��t@�$�8��Q}/�\'��ɵ�� ���aa�S��#�I�kl`���A�&���E��bY��
x�#�Dgǩ	�98+X�6=l>p�8�`�{�뾕3���m��R���AD�}˙��4)DP<Iy��S�W9n�����J�o0��4u�M�PC��|r��3l��br9�{I�	��·�~�Č����O�����HO�	TC�>y�o 2�X�����(|��W*/��T���/�����k2����J�T�=���m=[Hf�NйVX����a�9���	��"�]Y��o��{��UJ0%6C'�������>>z�S͇?x�fg�z����}�"�g~է�οd�;��>��( ���3��R�PC���~p�t����T�,9�^�}��B�x�Rp���.k-֐����:�m�;� �l?�600PI��d����_c���Ke�c뱜�����z�<@��[�d�`J�1Pʞ�cpG��8!A�+9��J�n-�a��g
��9g�jT<��U�_r Z���e�����+ފ�?�S�ey����X�|T}2g⦱Z���ӗ+�(tk�,�hc"��y��>��G�{Sxs��(�]4yc�;�>C��w�=P���p�93$RX_E�:r���+v����J!��wx_��آF���;X��D�/�����o�%U�4�,�v�����v��eņ7�x�QL�	��~\ �AP&��&gv�e��1��ێ�n*6�ԯ��������a��[��{w�<t�<ZnL}��|=y��Y�	~$��\�����+t"� 3X�;M�m��t;��7jS)y�v�k�S9q{-% �����g�}d�,���[��6��:P>]/�}X�P#f�V�4�ZL+X��w���� .�&�%�C�����W=UIp~�	�+k��N�I"ӆ��/˙ga)_YL���i�������s��u9A�Q�sG�7�s�at�{�&G&&�10������{��,@�����?�~��Fd�b��ẀPT�P3����{���շ�Ru�|��gzh2�,1rY5q"��M�t����Q&~�ʯ&��B���~���g�>�̇O��e}V�2'�YW�A�{���{�`ZI�F��ӂϢ��U����ؑ
�*�Ƣ�n^���~wh*��9��_��}���������o��ć�jnmF��:�D|��We
�D�P��w��:��*"�U��2��%���U�nc�MK�ح��^�q��I���uG� �^�hX+�a�������]E��$��<�6�R�ɫGz���3|���K������֯��`=]��mD���i�b%�ͩJe���rM��Q=ޅ�;Fc	M��kgO������QK��d�J�X/��x�P�D������T,/�*���%H�ϰS1?�wpC���c$��.Z5��F��k��7^0z�@��i��� �m�ZOH�s���<�do'H�8�{h
�+L���l"���UD��mp��w~�dT>O���}��΀�t%���附���Z{���Le����w�t��e��@3?S��U+KtG��jHY-���ihHb�c�Y�#�ذ#,�/i�v��و4�\ .�z�uE�
��q���T��v��i���}�q>���5Ųg�� ��Un쫎]��l$(ץ����:(�2q�.�?�D��	{7U�Yļjji^ș�i���é��s�)M����M�f�O��}`��܀r���~�p���#ܩS�_B�'�B.�:���:h���rz�P�3r}��Y��2��)��vJ��ЇVǹ�ꅺr/�Q��ca�o�ԙ�M4���ҝ���y�wʧ�f��֖�R���S�^�%<�
�"��v���}�T���q#�5���(�Gk��RB�ڪ���k�>�O�� ���f�	u������t����ky|@A�U>�IWe�5�b��JJ,�j]9�$�w�#�6��2J�Ŏ80�#ԋH��"���%�B�P���6���U�J9(d�˱�V����6�}�.7�MJw<�3c�I�9rKպ|FWz��wh�Ц���+�Ğ�i��
�toF��*�W�ڴ�@@�F&��aT-V�h�!(%��X9�lp���I��l��"�f��~3Z�UM��%4�(���:��N>=�h��{QA�Z�K�8���0�x�A[��d�(��K�>�Ğ�)�˛�t]�,԰��@�˝��~ܒ0�p��%gil�]C�Q1p�Ɇ�F�k��H"�g�%�!"��N���+�U����D߉U�^�yAk�}΁�z�dj���F~�O���\���!^u�'��0���^Ԓ�r�� g�8�9^UEq�D�r������
����K���<A��CWA4��ze 0Y��zw�fZ�
����[��c}�&�[JR�Ry#s���s��w����4��4�S��H�t�U����	87ŗ����c�'<�Yj?���o�;Eo�O@�P��z�Y����,q� nY�ǘ��ۯ�l���kM�(P߰�����d� ���u�K�]d��Ʉg`���I�2��u�m��O���r�py�t�#��ˇT�=T���~���Ь��?'�bϧ]��:�� W�)V���f�5�����cxfbe���)��Q���˩�Y�8&�a|��o\��2f4
|�,�	uǘg%f+M�[Z9#i �Qvy2��䦕b��:A�`?����ѝLW��(�K����`�>�����uos�,}�܊zHM�� rE��ruHN�2ٔ�n�y<��l"_��xd�S�����W��=�͎�@YC�ƨ>�wl(��<��Z����Z,���qA�����Pp[E�h9�[Y  �O�����fq���{$�����r��|G�U�R��z���p���a̕A�+u<yF�|�e�imoF��9�0W��]9v�'=�Szp�~�JG��e�X[���;��HFi0��C 5��.�$�	����a�<�?�~ �J�W�8t���SU�������H�W�<kӌH>V�� F��U�X'����qb��]��w#�z@��f5�����%���{��O��d�ꛆyL��ZD�u|����,'I��0�l�q,F�2Û�u ��&���kyR�ֲ�ˡ�2@j6s�r`��ﻻ�z���,a�4u�<�E��E����]��:R2:M���]]JN\��I�h���^�'�a}����ac*z���oMmq.�H73�j����dv�)l����?,p��k�o%;,͊��Sb����p�U�G��r��&~�Jl����G?�D���W0hvs��p�&�E#��rh.�%�g;�`�'^=�;�U1�����Ϩ�-Pz�7=� >�d��A��c|ZB��I�e`����uD�/�����JƼȜ�VO�U[`���	7B��Oϸ�^Y�*I��}w�޿����޴����&��>*�ޖ��;oI��+�UW{-L��`��D~~+�R�~D_է�	�'��E7���[�*�j�˧5=��R�q8��Sl�zOĄ�wk����5"c���y��-�#o���C>�|��|[�����[F��䅓��I��r�jߏ4�Ӿr=KB�8P���S�I�h"�4�����V�MU��c�;��3�/q�9��_ }|#�%���䷩�8���^���G�b$ac���rN��RZ��L`M����dUTx���֐��R���JQ�D&c/gtٷn/N<g�D�e�҈��{�Ti�wM�! ��GU��9V�ڪDU>#%#
��9�$�暛�D�XZ�����^P}PCWHw�n��Q��|����l�Vp�)���P���{d�!�'��y<R7Υ�E"m��]-����t�o>�]gt3_ڛX,�@
��������[�ڨ��(��(à6a ٝ߯���]e5[�"w�#&���OX�5Erͽ�C N�Y�g���]H�������Kɟ��+W� o{�hY��Qb]�a���/c�~����,s<4�1!�9){8	��YoE>r�n���T�����zeJB�p��#&ng뢈�v�q��]�����z�-��Sg��iBl�"�Q@)���gU��f$���}w_��Ŧ��(b��g�H�X�%���V���@�7��Jq�N������%A����u�2�F��+�+|`?���~ĿN�4��5 hb���(���^���h�Eߡ�\3�LS�3�|�?o�!z���h�H��.?���7AuwX�#NV�Y�,���|�0��	˪��Ikau��������#A��O�d�y�+,]S^]a�%y�&�)R2�z�r�(�#����Z� ���kA#��m��BC%�2�V��P/�X�t�l��O�G��sE�Xye���ҁ��Ȏ���$�i��Ώr=i�{'��v�Q#
7Y��:w�cѧ���8�=b��\^�-(um�std7uA1��d��t�MVD_�N+�Nq���k���XϖL�q�S�8�>�,:�cߥI��N��Q�
������+C}gT�|i1���|5@��D����:��#�w﹙z�!�*�*��`�H��x[��o]�|���l�
�+�!n�� �{B�|I��Q��@$S[h�fh[�ai�>���B���:���u[a�)���rh��L�6ϭ��9���i�u�7�+�G6j��B�
�+`���-2��W�����z���؁B���lp%R���>,L>�U��琹�윌��(hu�4��툶�ӕ>2bҁɯ��.�68f���>����gͯ�[۶�A	�]�ĐGk����\�p#u��Q�D? y�_g��ܖ?�����(@R�i�k�l
5��
�
c+����|Ŀw�P}jv#�U�7���m���/w7�q&W���M q g�Ip� �OcC��go��V���	cum-��$��K������8{.�F�����L�hϺmk�8X����چ�+Jq��|�O��D a��6Y=ۆd�?���	�.����
�����}��u�C�3�N�	����C�
y9p��þŎ$ܯ2��=��J�fK�di^����ƹ�c��� 	X��W�o,�X��ڝBF�N��K�x�|�X�<&��>!�_��+�b?�.~WZ��N\���6�ͬZ���`$�ѹ�X��4�(�X;�����B�`&��N;��^�acԡ.�Z&��������Z��T��dO��2�Iu��<��h�S۲ᡸC�-���g8q�M8��w���΃�0���+%�c�����e �V��vm�[9�����i������Q�����V�I��� �w�9�s���˃D�����������]�c����?���e�����c����dtO��:o#��	�z�������JQ8�'IGe꿙$v*.a�x����Z����D��:L�-+ϸ��ʹ�l�LPp)w�	{)ly'�/��C��"e���797�/�N�W(߰:��u@P��h^��@��]g�7�Đ�9ŭyQ|�f���sKM4M��w��t�n는��݌Y�-o��F�r��p��N�f���^����������7�8�J�IkcۂD��������"��}���-R���FCC(�$0���\�_6�*~'zs��n �/q��̣���?T~��E�UD�"�>Jt�?����L�4�nuT?~ ��Ð^���u_�Y�,��2:�uѦ6�+4 L�,�h��y���IM�Ҫ�w����]%���c�8�,�ןl�O~1r��e��L�方��{t���w�Ƿ��d7����X����8u�m[/Aҧ����1*g}���X��M��䳖�uq��H�}7j�/����Y͗�UE/h8|�0��&��l���eh%�����DϾ('3���������Y�u��1ߞ�h,e�����G�HN���#�gá�h'��� ]������h�Z8�Z2�飄�	����[�<jd�>���>����t
>�v_��U��:7�G��Q�o���c�����]N�R_�˼�r�:�Rfc�qaywM�կ��T��Jz�˖I���(�l��� ���%8�n]h�lli��5����A��;�?+�������O��m���VϬ<�N>�ݼn�{��-m��̞��o+��R����VA���WxP���f��cS
qu����8��U�,��^�4�f�x� �-N���������\��[�@��L��i�M���V�B\�no�"c}!k���5^H�ɪ� �F��-8K���>J�W����y��M�����Erݷ	H�|���Co�}�rK[�����(*��#�dAh���s-+�&�F4�X�y��NB5Px
�Dq�'"��?�Gb��L�#����8����΂�J��q�E��� Avj議7xȁ�i�C���a��l���n���g<������#�� �7�%*�0ͽ�[CnKo�+Ă�8�&i��>��M�)�,��m{�-�,��2�$�	&g.�i�0������2&�o6ik(�L���E��d�u����ε�ӑ
��[�<x����s��k��G��cK-X�W��[m�=�2����9P\-�V�� ��Zk��Ҷ�ǯQ��zﰱ���s�q}̡�A�l�JɻV:��0^��X�ndO��6�c�n�1|���e�t$*8��r3!��߲���E{F�l�k#��P{z�:~cN�晙��y4SQ�[I�1�Y�R�m7mo��u�u�RvI�n�U������G7XO��S�B {6�4�L@���nM��m�|���4%Ӗ��h&�4��m��3�.���de���VV{��	�(8���xV.p�")�(�h��e<wX�i���~Y�#8��N�y=86�E����n|�a����������L9��f�I�O_9�
dr��#u��Ļh�����e]r�Gh���2H�G�F���+��!�T��%c�q��ضy�R>�|tۤڗ�v� qX}�4����t����έq��m72S�0WVz�&S��E���2Qܒm�TZ�%l��I���˔�۹}��&e�����d�̒���B��*3�]@��=M!�mK��Ih��qsq#��^�6�h��� R���Q?��i._i��f�}Et@����A ����78C��;�V�b�'��a����`]�*l�9�6�^���k~vP��X��Y�r!N3|��4hMc�̰"M}E�Aػ;b�.���<܉$���x���7�7J�s��n�r�����U8�Z�捣5P��2�V�p�k��N|��N}�J����L��Z�X���6�B������C}���䙊��k�\m~�%O�ȅrO�DʉԆ�;nq������ۍ}�e�m���xb�Ci��`6^��rJ��9y�������,�4��*��ݦ+�հ>���h����/�r�7'a���[	�@�_� {����V1�ݦ�H��/�6���4��o����Fz��j�K[��&���]�#oa�u�����_L�)ڋ�ℨ�������և
n���8���>���!��;�!�嗪Dwo��A����ӷ��b�n����FC2"��t�9���a�0�׼58gZ眈~~�Eҙ3��Zä�I������qI�:,x��>����f�J��>�<7ѓ�Z| 0`$k0؄�˥ �'W���"��+���\S˅g�Fr�-5$��%��#������6f��A���?{�[��e;�Q��0��Z1+�Q�ޭ5x��[�(.z�I'�I#*���*$%ɉ�v�\[}��l��y,$��8�?4v�O&ƽ�p�d�Q�P\�m!#&�T#���	y5�T��.S�Q�0��� 6�E��V�2�?����d~�~��Ȱ��jz����ǯ�XG;z�=z����/�|����qr�S�KTe�8y�����r��l�|�	��:�������M&UU�֐_��3u�U�yY���x�I}ai���h��r���9C٫g(D�m���^��(�u g��y�G#�`�a�S���1^��ȣ�o����8�/��B����2��}^��ϰ��eq�<�����w{���ԴG���=#27�:�57i�v�[/��U��r���з3�׶��Z^��8�[i�U˝��_O�Z��EZ�̭�1Z�Ü:����ۼ����Z
�{��&Q݇����:0f`��X�g�6=W|kr��Dq�Q�^H��\��_��Q��m[U�'���	�O,�Or7�c�����,���/�(:9��ӗ����e�X9�.Y������V
�ܠ�{�wN?\m�Z�w�yp��='9��\��Δ"�_�H^���J�o���fn�61�|].�R���'���n���*KH�¼��jjk�=8��=����S!�k��-[
o35�����}�͠D��ʉ2:ͳ��N�S�N�1����U!x�ݪB��Ҧtc��`��ŧo��A��R^7eۜF>)�u����cKo�zQ�2��P��P� ^N������}�_v���c�[�,�����y�W֚�|iWr�ջ��3޽"'3��KQnS+V����z��J���\�AF��L�٭�l�@.l����ܶ�H/�z�k�loT�X}(D(��#o���Z�~!.��]}���zG�M���|k(������{�����Q��6fd+��3�$Q�����݃$�d��dKЂ"�A��C���c��BE=#[\)12�e.�g����֝;u7Ζo4�`Q�W@)�}���,��u�'q�#��a��[M�3�zȡ(+�6���%�V��Vx;��x��dϠ���o��P���a�.l���?��ۗ.ig	�}g�8kx~&���t�%��֫��lg?�:���jK �^߾�5���r�������b�
�Q@7�N�R��=�
Q,���;��������<�l��ߊ���W��P�,��C����ɓ���&��i�C5^�m��l;�j�C;	fj���@o�'|����2��Zmn��C�H �W���o�$O�sF|��������-1֨�o_�X<f4S�ߡb��ײ�!A���9��S��rԘ��zD$��]��i,��z�4���f����C��Ed/�k�>�-�B2�P�}�Fr��Rm9�x�J��1yW���o�C�J��MѣqK��u�cjPs9'��!\,��_]L�kÃ5��iǾ�@A��&�^kI#r�r���9I��S� �]
���P�j�Y���rtG�.����h�y��Iy����㓇IB�Z;T���S?���BQ�h��h6� ����5qn}�6O����"�;��T٣΀�ɸ/����@���^К�4��yﺏ��ٓ����mL��<����9%�
;;,v����G�!}۽-�L颅��W�/ |�Q�N-�Y���dה��t#��KX�'V.)�c�{�Wdz���%KyJ[���Akcj�J������i������)2�H6��]>��m��${���(��H+̠���Fc�r/s�xIX��L�����ְ�b��D��^�JAf��&�
��������*�O	ޚۿ�+h�4G�Z������i:�6u7��/���M70R2����(p�����B^(�S�q�k��`���Xu q�h��M�/KZ��Q�WG��2��&s�'+�k�ڄ�w�2o���@�/C�����m#�֌��&F�Xi��[���`��fa�um���܅���08:��.?�Z��6L��W@!�j�@����Nd���#�iHh������]��'��@��M�������D1C'k;,�m7����'@<>	&�d}�=^(�U´��"���p�
��:��	�tW[x�z3Y���ff ��PZ⡤��D�B�w��� I��"�j�0�����dݹ:{��:j���������I��_�Mӛy�R|��3t`��X�91<⇳' ����g]00<�Nl�d'��mp���r��?��%乙<�Tzf�๭�V�J9�={>������ ��y'O�j9W�[Şw�������\%A/>u��?�vǻqE�v�Pd��HBWu����YB1t&���]�f/OWcy�ipO�|+��ig��\��"c(-�h/8D�#qʖk1��R���P�HI���u�%�%��!��
��{���)����4��z
<W���f�ڻ��օ�*ۉ��W���7�ꚬ�
��<��'u��k"6w��5��nqg3x������$��*�~�%ry�v2יWq`���څ#�8��7%�U���N�J��3�Y��uy�7kA�#\�R���'꺏���u'+�ߨU6�p�^s�V�E9�L�?�L�"��:x(z���g_�N�<ߛ���'ɿg^�� ��;�'s�n$�W�˽Q��@�$��t�'/�C#��+�k h�=��FsS�k�sAjjf����r]�Кᇠ@�˓Vw�f���z؝i}`��p���ډ8L�NQ-i���,7 \�D�[2Y;tA!�/�4>SV��=h�}®�e��׀�O�-��������w�p ������V��O�[j�L�˄�+����od��F����*�
"o1w��b0�tㅶ���w�/�'�qY~S1q;�u��\ʬ���9��}��+
W���U�/����J�L2�^]�?P����V�Q;��-z��ܲ{�ѹ:���2X�i�
t6���1B�����K���9�}b����%Wj6xw|��m������,�|9Kg�Q�I���4�Q�]�y{ΐ39{�CM�����2�fCґ�d�;dgP�|�B�H�!-<������g���45i�l��H�nri������׀g1U0i��&��N�;��6�&C)�]�ֵ'K��n�Љ�)�S��T�c"&>��|�@�qe�,Aj�kC��/_fk���6oT�9����M�A����RT�_�?xvLxӸ_���hs��ݻE�������T+�Z'߾v�|����Wu�2N�ޓ�5+�a��zծ�lb��G|L �;�xEvǳ�n�`�0l�ibD�o�{)w�`��c~���kd���t����5�y���D��)�g�����[�|�j��`_��D��MK{���eV�H#Y�s��.�}`���.�b%F-����h��� ��Y��('�p	��T�i��� ���@%�>��~٦�����y܊�r�r�N]t���0Hcqv���߈ͦ�E�^,��SR�xW�Q��o�xn��9�c�tA��lQ
�2)��=B�1��B�|Z��f��\~{D�we_��b���XK�ڴD��ֿW>]���>1y��_��2Z�˚����4˷�'������QC�������I��"��ٻ�}�	�>jy�ڟv��ǽz�7��<@]\�O�KW?
��%+<QN�V柚�1:)l��7����ӶO�Y8��,ᩎA���	5'm��ƾ�ׯ�t>������ӭ��Ԋ)�2�����z�Pk>�^�ͨҞ��\Z���ȔOQ��۾kw��$" 0�)�|f$^*�7t.����z�A�Hd�����m4�X߯x�TL���!��I��|�^2��p�����%��vu)x$�|ɦz^���{�\��N��@�u�t�o�������*�"��'U��9t ��5�븷�)�@�@Al��	�mओ���}���*U�5����N�g�Cwl��ulZ
I�c�Dc�(;%�N������i����"��JX����L�@�<�@Z;us�[���E6C �2kq����$+�(�ߠӓ�gH�1���"Xk�MuN�p�&�y��äD?��.'�93�x��)�Z�WnL�M�=wO{}dtz ��d!�y��Fy�r�w�̬��9����E�V���`&&k�p$�c��=�eN�0c�\��s�v��"����/#.~l�ư�� m��B?�3�4k��ٵW���@�x;��8u��ۆA�9XA�W�n��C+�t���>��z��bw3Q��w�a��fQ����zd4|%�7�Cg-�iB_�n��Y�cd b�2�=7k��y����b���AjՈ����T��5�Ơ<��|C�!gNV��5qWï8�s������A�!R�cz3)�o�C�B�KX0owN�(��×��T��{�AK�Åsg����������VI��)#&�V��Z6�[�u�KB!N�i`E1Ndj�$��p��<8w7���Ѳ�^�c~�b�=�WB_]�'���KJ:��.h��ɘi�<���^0<k2��$	Q8u8�϶J��*��|�B����ň�fö��*�����	�/_>��ج*�兔�xa����������7)*�o4p-�|xȱm�����d����H"����@c�u���1��~�x�haXDd�(tZS�>X�?�Zƞ5V|�.:��Gւ�@N��`��p���E��8�ۓ��$�=�ȁ7�q���V��R��(�BK-���C��o~�6Ԝ5$빼����\�0�	9xt�}}�u�u��A%���L���	,�<*�_1�ѽ��hCW�>�<�@���B�T�=��S�-�9J|�MW���ct�OZ��m��������ʒ��>�l�k3/��t���M.�FJ��#�4��
=Q����-����:�Al���W�h�@,�l��aZ�����ƃIX��Sj"i\�NS��%O�rDߛ1�5	뼳 �ZC9�4<4z���r}�ū悎�B>��� �$�a�>E�˴�ٝ&�IPeiyR3au�C6���w�=m?'�8	0��|����͌�R(��RSjQ����vJ"ynz�Z��ۜ���CC~���-��%��C���-ȸ(�P��l�ffGDP��UMɔ���4
A�d�
W�4s���Ӎ���@�*.G�h� 4�T/@\�jX��vnz����C��U�S#��>þ��Q;�j��> �V�mW�aF������7��uG���3���B~�b{�Oh3ӣ?��r�DUD8=
j�倴)+�$Z��w��c�zC�8�aF�'��R���r=wNO:B���E����G�z� G|j��i�{Zˬv�rQ�N���nH	���w36��Os	���Qj6E���	*��i�sj�F�F��{Mߤt?V�#-����Vu~LEX!�]-����w/Fʾ�$�t�bR%��l����)�w0���	�[�e�F`S��C�Jtα,K�S��B6���fJ�����_�TF[_%XX�!���>:z�GlE"P-�	��c�ݥ�v������?�� ˢ�R{���MM�]2Q^�G5t�i !�j�f�d�1 ��5-�6��������֪��zX�Ȍt��#���v2�G�x��R�8�b>`����Tp�C��gdqs#���%�M�����ʆ�c[��F�MoK!�[(��
T���H�����o�&6�1�*}�8��b�pV�q��Mk�V X�_���U��:��F@�~~�cԛ�����8�m!B��x�N�%��I�ii�Ii�h����1��eF�~(�h����hϤ�W;5Ly�E�􈩻4$�9��M��hK=E�NSuAH����-]�α�~'�qx�U�A����t�{�!�)��R�6�x���V�ӌ��-NSZ�Q����ٟ5btN�o�pČi6�gb D{�����<��Ԗ����I�53�9�`��lAk� ���7���@�(GI�3����O@��C`Z<T�r2�,>��$�<`a��d�h����K�]1�*�C\�����*ņW{S\� LGv�Ak��.�2`Ā��~pO�$�,O�ʄ�A�GdXyعk�Pn�܀�#]�9���٢'5�'��6��	|B;$J�t�b˺��,T���#,ĞL�.�*w�P?j��DQ8�v�O���3ɋ��t�
5������x)i���~&�&G�N�0M�z�z=���Q ��:�"TC�9P)��������c�C�T�z��~�����T=\
��Wݲn�:J6��q'�mZh ���{Z��Gߡ���ꈯP��#�S��4�ۥV%�@ o��yO�qxZU`j0���h['eX��+=v-��zo���b�P5�͈��Ix�ă�R��'Fr��\��V>�	���ǎ��5�|ݒִ�"q8�43�0�G^g�$q�zq�|��}G��>����Ӎh�����4�J��P˂��K �>��n!.Ƒ����i�L̟��#�3䃮ټY��C"�D`��!NQ�)������Ѣ$5�HQr��ߟ�(}O��NZ`��]��|t����1Ϩ(��n�~�jA�0ҫ�2� �U��� }y�G�&�;�#6�8	(�[�ux�+)�T�>�$�+7U�d/P�N���>���a���V`DE����ݼ ���Bph���z~����3��U�1,�w��S���~�<S�~�O�#5�m���N
dm�����	4�獀n$�5u4�tt�Rz�5�S5�k|��&��ϖ$1R�O%e�<��D�G�vᗦ_<2_5w�#�g ��ϴR��̻�,R'��,�Z��d��J��H�����pqf$�7�(�&�X�^D�m:zCX�γ3�(Q��(�l�/i3�~��ZS1-E�V8P���r���$��BտOwo:l�D�`�R�ʡ|�Ł�T�1���ׅh9��E��e���]5�ħ#�r�O��{S�v)|�RWs��_����	/��Л~k�����u@���:�UCۈn[�Ղ��F��ʪ.4JGX̩ԥ�d�+��9�h�3�R�hA�vSN�eΎ`l�ڭC��N�tCO5��Ε"�=@ԤE���7?��H ���k���!p�x��Z	�%�7/�6e[
gīU}u���?�Y5���R�Ju����c|�*-�?�g�+�'��R����Y�ow/�-�~�Ԑ�7�X9��q˥E��XaU��0�J{n�3���t?��'oI�ݖf=���Ԫv�%(*��Wx^��z���ϓ�tnI����įCP�ҡUU����2��)Yaxd�_A��e�\��Q�	/>`���М}aKMհv�!i�e`��#(a�' ���+�U�I�)�a_L氚��Y/܍���?�z�`����x�0v��ǰim���ds�\[ �SL#*}ӱ9m'��x��ؤ���@u�OZ�n�����s�_ֺZ�땽=9���Bn�������+�FA�궝�٭�{��6ջ4�I�8�Rd�u
 �Aٽ�� �AF�5�Yt�>���z�R?b�y�\D��z�  ���ڧ?��H�K�H�٩�}~K�4�|B�O�}� u	�_yC�M��"(Nc��о����:FZ�����߹�A�Z�E��[�%J������C�Z1��!�� ʸ�Ȕ��'�#����.L�%���{a��nAǳZ�٧����4c�@�%�.6&+�} �Z����h���"����_H��%�x���2bRE�&Tӭ��#�3lL�pq�D)[���n|�m�ן*���XR �}���=��s��R:p�^^����̽���p�{A�F��n�'৬2`�����B��i�҃��y�׽ �����Rb�D	�Rŝ��SuKǕMf��"���I|=��%X�]�L���İ�т<�ه��c��(6�"��.�ߡN���\�cX�MJ��B��55B�d\�y�a��WZ(��{�z� �a1���9��U?t8��=G�xk��ZG�:�X�.T���r��KkR>C�4)]ТA�P�u�4�9i��i�����Ǫ�5�15�`5�g8P��
v0�8T�]@�#�����3i�3�/K���:��PLEE���ao�=;��/> U?$ט�d���j�v����H���K��gl�]�h�ŶwYaVq��bү���Q��/�Ɯ,뒘F�D�Q�_
V�%���W"dwcJ�Ӌ��$\�߽"8uK��bPū�1W"375V�"�VA$L-�1(�[ɢ���r^舻j�4�ܗ����͍9�7����\Tt�\��FU��W��̝�s.�3�w1 �z���J5�W��L��W߶$Y'���{�C���)�^x��W������A?~����)� 'Ѕ�)��Bω�K�j�qp����tD�0NiÑ~��^�O���w�G���m�Ì�R�~�D��S����ғ�ɛ��f��oA��n�&��9ո�k�Q�<��o��¬��{i��q�*��H3�EI�$!J)[�����Y�K�	�s�2�`{/����
#}J3�83rM_Z's���HJD;k��HH���HQ���t�!A���ם��C�g(�F��>���S��Ӽ-iZ�pm���� ����@(��MU�����]�����)��^�e�"��]l+:�u���.�{Z�P$���Tl������aM]��hZ[m��� 2���Њb+�2*�(c�A�[��(SdT1PQ�BPQ�QE�0	B ��a��O����������}�+�Yg�5|�g���I��?�m���4F>%��ܜH��=�Bh;�ejmY}����7/��O�[q�됪��
n�lP�ԉS��m�h��ڛ]�7w�dk��׽|\貴�Yd��U�@���-j��C�e⠅�й_u�|28�|y��S�}s2���smk���e��:�rvHTy��g=�/��(�ʬ��OŊ.�kyw�ls<ӫ��/m͇c�Hq�j�EG�Z���lֽ2'��o� (;:b�� k�p��@�vߏ9�#G��rx�6��	=l�B�'��'aS����h������8�s���M��`hQ��J6�J�J)�1��l�D��9�c�qv�L�����������ϭ�/v�/�r>��i����9�F���bi��%�zƙi	�������f�����,fgm��F{4�[�$����wD��ԭ-j�Vv|��\��ݦ��.WC[���y\��[��_p�*߼��ě-S�����ܤJդ-�E[��Dq�X>����L�;�ې��W�<N� ��U�yZeg�ޕC�[�
����T̏���7��h�f?3-|��@�~뒔v���L����e�s��=��1�{J�Y��U��AZ�OK`��0�i��EO^�������l_�4���ͻ��E
:m����s'ֆ������ZG�$fc����O}��{y1)\�%��{0|��&�`�y��Wɜ��6�:�z���d�o�8s��0k�k2��x��s�ܵ����6-Ky� ;4SS&���,�^殝/L�����{�%jߩ-�a�u:��ȑm�ʛ♃>���9���������^%����T.���,¿O0�;���Ж��33EPĞ柯z<?�2�=s���v�Ѱ��<U��"��Q*tXlp�+۫��4?�!D�[�6�Ŗ**�}_w��۝��RO�ދ�i~I?d�Ie��~v[2כ:��O��i{-�Ś���}i����u��p �_כk�����O=����/�&hs�ν���}jA��p��@Q�v~j��h�1d(9�;�nBU[��T���nm9��7��`���#�ˬ��]��׾�������pq�Hv�ýYy�����	�l�W.�E�8;cWMҽ�of�w	9{~�DŰDf��~r�~��!��y�����u	�Ԥo�b�;͹{�_�7r��{ʾ.����V��Z�t���]��u]4�^q�`70λ�og]_tF������Ӆ<��;�.�m[5�8޽'ӣ��2���o�.O�jf�0P��)Ӎ���C��'�L�~j(k�}�}�77�:ER���~���;�s�����ǜTr䷩��F\J�T�ޮ�����-yS3@���+cͮ��S�N�8�q	���5{�G�Ή�,J���4�j�T�v�"��U���xV ��N
\���R��&l(��Lz�hUJ��#���;��O�+�3U��Q��K�yX�|���!-�
�ڱ�'jS�g9���>�{��̥v��q�J����Ɨ8�֮��`���_u��d��>���gpx��+���\�l٫޷��dC��EL��5������g�n�����/��uM��ph,�S���+o�B����qM���������vA�o�dR��K��)���;�|���t?Ns)���p���;.<��z/��i.{�+�}y;�7���~����<�bx�^�H���r]����.e!����Z��4�8�^�tk�I��r��v����mZ��z�K�ք�}ג<���潡Nm/G��-ͷ��o	���r��hΖr�K>o�s��%�ʉ��-�Z�g��l��q�~�K��ŭ6���s���Gj؄����)I���Ι����)9�)<14��z���ӷ��}i����]y����H�H`^H_E��D[H_�&
�1���Ɉ��iZ�;��o��~%v#ʚ�$� Mя�2����oP��m���K��\���/�~��˥�w/��qBO,P��d��OU��|;���Ҕ/��������Wj�7�Y��/���՗W_^}y��՗W_^}y��՗W_^}y��՗W��yu�w.dK!GdJMA�KS��{�2O���m��K���.�k�����?=PY~�ǻ������!L�����wk�����k����oB~:�����L���Y�~A�����I�Vao˴�̷Y)�)m`�]��qj����}y�˛_����7�����/o�?��?���&?�3��x�3��?z1��]�$��#����X�/o�������k>3OE)�-z"���g�������շc���|֧zr�����8E|�Siy�E�vI ��	������2�DԾI\JO�<���k9t�,y�����p�h���s���Ѓ?�Q�"��C�R"�PI�\6�(�<"�=���g��ѣס��m����z��OD��&+?�<5'���[Lb���;i��Į[HE7�3{S�<:�^���i��m޼9+��f�\��Ku�&Bۜ����N�/�8�$C<xO	]�?���"7��\��g%2�Se��hk2�������n"��ۻnjj�[�siR�C޶�:2N�Nh�:�?��c����+n�W��}p�$�������������Θ�����T/
]7O����p�4鈕���F&��@�/��Z�-K7K�}��.iߖ��Hj �t�M��;c�*X�l�~�\S���ay\$���br���w�����c�}"�1A���8�����pKb�[�1�R��M���J�}��t����oi$jW���g�E˒���^��[D��Ik�=������AcHl��U�Ħ![E�hS���h���2�g��y�s�Qe]�(hI�1�1�q?7���W�g�Æ�>��W�|��pV���^!�m���yMϠ��իW���5�˰�+z����n&,>D���FE2�M�pd	s��1s>���<���tK�pw�@ø����4C^[�*�~ല� ��Pu��}������"�-5 D+w�6T���X9�����ACiP���;88l9ED7�w9,[�E��E��2\�Y�-�sr�ख़,~�DTم[��[0V=K���z?`�}u������-*��*�ΰ�.Y�c�+�M���R����g���g��/��u�~P�囦�2D�	=��,�4%x#��f�<�W�5�K�|�2�y�񨻅��s��!�_�f���A�`�/iPAN�^��ж���$B~��P�/o��L �B�b�m�&��q[kk�E�. �,y%z��U<Wy}�3d��eFKK�VQQ��	�����p���_^0��C:�W�V��߫��<�E �Й�}3)��?/ ���\ ��2m�֣p��D�U��aq%Ae���8����!e���A)nO��2÷~z�����������/�C�e�9ro���x;��t�ޞ�@�{���M�Y,��k��̹�*/J%l����D�����nT�Bui�Hӂ��|Ցp;&���KH% ����ew�SN�*����-(��!��K��Nu���.#c
p�uIII�	i���pDn;�&�Zl�i�71�NH�W�~���l HЍՓil�v))/��B�4���(�[JDK[\���m�oVf���3_��	8 �ն����7�.�$PR�����ϻu+���D�)�%�
�]�?6��;*�T�\��>��!@�CDn)-����@0����gW�^m*��,�#h)����p��❽3sD����Ÿ61+�|�/%�8�ŏ�E�QT�B�܎)� H�{co�-�%�����'r��3X�O���(77^� +��řC���g?��&�q��DW��g@��h�P9�)�-3v{�;�mZ��v{5튗�ci���UQe�D�7^ěj��ڝ���`V���Mgl�WDk��R�j�cuzL1,�+KO��j��}R��g��sZ���ۏ�22�#
5�!�w)� en(R��f��Гu�?��x{-~�?m,�v�l���b���p����ɪ�ʁ_��|�r|%���&�}b;����:X�ܮ��y'h�_�݉���yB�(�����񴰘G&6�+���,�!B`c$r��Q�W��Zʒ�y �bD���V��+?��͡������7),) Ȋ�*{	h?4��$���o�=+���޶!�o��8j��k�!��W���S�� �} ��[��m�����
kjfP����x�X�;��Yb;����I/@$���.^�i�A)��scN����̘9������"D�_���9���/�-�R�[��r]l +#rǵ�^5)�!�V�,_y	�L�������N��>��ծ����;�-h=�}�X�R��x�Xg@4Ʉ�N���X��!��*��M���DsCh�^�Kܜy�Z	r�$�4J����B�22vh�g����U�"Q;��X%��5��AU�e�9)�D�� ��k >�����z�F�N��u0��B;���� �ʄӕqT  ˣ�v�yg���"�Qɋ�:��ٔ�Q�E��c�hY3;�n~�F�^�<9��K��4��u��E+�5�5�u�����)p�d�M�)��׳�3��Aa��W���5���H=7������4�؝�O��>}*SUQI�D��a��iYY��tT⨶��g�H���jK"����f�0��P�ξl�΍k���y@d�|�ȉ�_���IM��=k�H�r,��	<:�<�,9{$"}S�����+-a�6���Y`�^���X���
k^0�x��#��0�1�����C
I�~,�l�%�
���n��	E��Ak��1Z� g�.�����PbČD�4%����G��NĮ}{�X�����y��%�E|N�l%�"�)���Tu��ح�|�O��bQ���Ot������������c�&��?$���[��XX�D �WOں������?� ���YS��3*+�EK��� *+1**�sx�$���&Q+��2�$�W���i�풱���ʽ�!���^�F)�����m�P��u��G�$�"#��+��(���BX�$��>�z�{� K�� ����	�BV�j��ت� x�2��#@Q�o����`e����xG�:�Y�Jeü��	է�#x[K�6�.�>S��X��m��$���E��%$�猱�����ߟY�C8���ХK9|F�j�@~˽�$,
;������l�M|W׿�.�������&�A}����زjϞ��2���p�a}i=	c��o�v��>�X�ϙ7I��Ą�QE�٩��k1���oD�w$�͵Khx�Oi?��ϟ�8yYY��;�x�}#3p}�J�tn}X�k�����п��HƺW�Q�_��%���)�������f:���)I���������r���LE�!Z){��p�X�_�r`)��4T4�������������K�u�@9�U�dm�(�`��i��4RY ��3ǛR~�ʙ�����ދ�p���x�;�)3��,�KU���@`#
��ƅ"��}a��^��˭_Q��3g΍�V����~UT�&̰�> �q&����7n���,o�Q�o�3p(ח��Z�c,�E�^��x�ňr b��m��>h��]	����0k �V����y.�?6���޵�n��૓����y������0�	r�.,�Z^^�.��������l�v��/�����	��e�a��v���(h�\%o��9ɧz�����(���tJYRkZ�1H��j������9 $JPe?pL�M�@�_@�\� ��6[;9���k
�D�Q���3snu�����%b#i��c|�q�G� f�N���sXfN[�~���B�� �JtV���|N��q�?9�xɥ�˨�p�v���'�@ǟ"��V����ʃ�1��· $H���k�5�U�s�>�l��Ǌ�8B�K�^z!%�!vV���BA�#h�^�i:���s��5Jr��_�e�X��!E�w�Ct��t���:��1]x'����8w�1>�:r
m�*��x��/�BK���KIl0M~��f���	+�x��g	��o�S����	cbtS�'_+�!��$^i#3fsH�;���j��b5J��Ή���"�C(|��fl��׏�:�DԠ�?>M����Ud�U�!>G�'3�x2,�� 2��!S������W��Y�X�V��X*�9!�)[p��ݡ�i�SB�YgB��8����WCͯ|��ٳ�V;��2�xGGo���ԑi���d��J?R�� ����2s�B/Y��s����y�JW�X�?x1'M�T!$�m� ߬A��O���y��R�f���ި!���z���Q�C*�i�A������'�S-}m}�"��B��=���<U��o�
���ȡ ��Y�F���h�x�3/4�g'�Xi)(SF+�F�K�ĩ��8����  �`���Ϗ=��%�{}�@~;-X��������
iT���2��]��cn.䭓��ݲ�-PMޢ Ʃb��Os�i��
C��|���\& (���6�*r�m�Q讁�:-���9id��"����w� ���X�7ۇ��كB�1%�J"�g��R��:	�yj�T�Yy �]��
��$��	5�9���J�1Cyk��;�y�o"�M��Ӵ�p�]d��9���O�рG�'I8�I�-��A�J�`2���ƣ���۱�L+�?��t������)۴�u?GE�q@r�¡0F�K��y0�"<ŭ �13�ʼ��k�Sf���p���b�#+q��r�� TZ�f�O��v� ���3sn��\�Y� �.����s���[PxӮc�\j���RԐxPN��Z�k 2uE�\��v�VE�vKu(6�z:��F'���L}�WD���l�Ӝ;Ϙ8�,��{���
�����o���ݪ Oh�u�^�n��O�'x��}NA�~ϤAM��7��� 8Ib8-{Թ�b��c�SE2"9	-�=p��
_
�/��4���-���E~�\�Y&xdV����"
Et9��^��Y�e�u*��6�Z�	������j�vN�0J���g=<F���kP��b;�LM2&F�C/�����	��6�D��{D$T�
:��#�i�s��Ȣ a[�wk-��?c[�#�5�+�!q0��������$����o��.2&����?\�z�汧��~�ƣ	��b�K�H!@%��$3�>&�X��fnȼ���IǍ���ޭ+�k'���S�ⱄЩv���HF!(J}�GǾV�ZM��>x�ђ��;��~�Qil��1,|�����`$�u�K򮙹�'��J�?∝�{$I킶m���`����#wza��~�}�&	�����W�q�S8�j�8�V��S=�y�vd�|�d�$2��̢�R]�cP(u��|����'�q�c��g\uYcӳ!��)����Og�+n�ZT�_v6�%M��Х��Qb�L�~E<�au��ߊU99�!95ɪ���a���8��m��V���E��S���� ���I�{�ә���8�>�$���E;h���a�OTYW�ObBMI�\&*��u ���f���\x*]�i�#ր�YV|^��-3�geI�&�?|���'�>�Ǌۮ-E-Cb,�;��]\\��&�S�r9q�[��Y=�:ۊ���Lԧ#g��d,�4X\	8qA�TTY������qMd޻Ȯ��
Z��dyRR��2d°�Ȅ_h?}����c��q¬��A�"g$^i6�
��K'��(��ޑ�)�����|,	�@��kwm)��nP`2233�P{;�ǣ/�C���uH��n���TUUec礈Z��2���yYء��$1?��YL����U����z�V�Dab:�^�#\¹4��be�m���R��@�]��(hF��JD[ʔҕ&�h�ÒQeC�);Q�$�����,�9uD�u�f̃:������� ���w�7oN[�0@l��������H��]sXy)��XZ'�𡶟.�����T��N����J�*��?{H�v8��^�N�"��=��h�>�F<~sk�ʂ-ʞ�/^���ʚ��W.�
~)�|Xgf?,�)���e�8� ��8<!��g��1��̊ �1
%�;�
�xC�U{4��?��Ђo�9�Og���C(NwJ��#Gޅ\dp+��/̜l�-Z ���J�6���a��d�� 3,,��1��5і���o���'�Cv�梠��?����$��Ц#x[���Y@ouT��_���\�R �מW�,ʘ�m�|�Q=�\ҿ�T��$/D���,�u�4��\g;��Q(��)�QjE�K��W���tf�%F���_e���us|�}x�����Xm����W��b��J򠏘�4Xx�ر�_Ѵl$������D�S���Ř�kʴ?,(�\G����i�F�㝌����L�<ʚ��k��dD�u_����Z�%d���c�Eր. �a������ أo�|\ǌ�b��G�Nt6���b����ֿ:ˌ�}��#|ׄ}�L���<ب���t�/� z�i�m�F���~0܈����z-w�\N����T�{ǧg?wN%�1���J-?Q�`�G�N���FK�����7b<�P�M�A������^��\�C객]���*�v &�_[#ʺ��z�����1q�ݻwU��ad�}�+�qX�}�I<EGIA�$u~��װ��&(U�	�<�H<��_�>����3/`	�>Iq���_����3��[3!8���C!�U��#]e	�	UR��U��nD~	q~)��
n{��N l_���u�9�(��x���K��wiM���o a����T�5�+��P��}��	V�-GIk�툫z> �P�z媉�/��%�!�-(�� 0t
�����GQ���O�+4�Ϫ�A�C�a~��몪*E4w���е CE���o�I��!4���:+�� 0�~��d��(c�9�&%ň�-��Z~��1���G�t��m׃��a7�N{8%�5��R*\%�?��+���@�}9�gb61c* �x�*/F�$Q]doŸ6���ǎ
+��̭��:��\��:���^�ԾȐ��U�g_8�
*��:2��AČˎ+I<*��Z�"'��/j�֏���B�2���(n�Zch�|�*��K�x���D�R��#��4M�d�#��kkʄ��b���_`h}cu�� )�߫����sEd1<�W���OAg��v#�Lau����q�?�@Kv���i�-���)��ege��[�U�`������6��<m� vSq��֋oUP$��lK�ϓf���V��Ȓ��#sss���A�[�7��#���/,�ӳ< {_4�������Eʭ1e0V7�[�)]�=�@��rUh�.�:�!�Vy�wK��D�g8����̜3+��-pe����`����� �A����QQFEM$%�`'��<��'���u�D��m�W��}�0�mѐ�����i�ԅ��`�%�W%u�̐~V|B�[f���I`��8��\�h�H�[�:L5=-Pd9 J�=�,���`pʥz8��[�>LV"BO;:NI;�����:!��,u$Z�-C��}���+%JXt� �y��2(��Q�є�h��B�R�1R��須��׮���}�ە���3ێ�I����3 ��� ��Գ�
��<Q:���kx�K�;s�LinhJ�[GJ<xp���쟌�0�a7�Xz 	=B�9�=�픒Č6u����Ð:R�����'"t��[M��
ނ �L��K4�"g�XsΙ�Z0��p�m%�R&)wլ�Os�5c�j�>R&w1.�F$P<��_[S�䟢��yk���>#����~=%7w_��O�ʡ�]y�>F"M���a�T^|�>��8�RH�~5/3++�ִ���uS�$��`��)��1�:�E���?2+l��Șx����3�܀�������bј9��()�߄1�9fD���v !�׹�	C^�n�;4��m��)�����n��t\��1>EdV�����P���=߇!{�G�������.'Ģ�W�t�s!S�Q
����cd{n=�Sy��Ր3��uT���`'����������D�y�_�CJߋ��?��P{�]�*�Py�L�t܅'��@}qR�����Z�i>�r��;c+�G���\2�$a#N�G	���`���9-�y,��/�1��v�'�e�*��
�h`�X)�����</+�����Q����>ϒ��l���g�����!?�n�٧V83� �'���W(~��Z�s�`d�u�A^�
���,>گ>B�Tr$�L+��~)<R�GYp۹AAA�(r��E�j`����?�T1��k��[�Mf�5�3����;��A��.)�ּgfК�P�Y����Ϡ�SYrvY�E��s-6vo���vx�絎6���T7>��^��Z��{&s<�c>��f>�y�PUEE��;��(��xVC��:RhU_P0A��������$⃨G������.�)#.B��:�Q^�l�
��c����9`	��cS�2?e�m*K"������`0�>�?��:��w Eb1f�*<Ƞ%�s*B͖�2�]�09�|���
l[�X�q��}�����^�z�F�t1<H&� i(:�������E��P�4�S����z�f��)N�{q閂�לɵ�.���*�;����J��Sr��0Q'�r�cA�bG VsQG���
����L�#�ŷ=H��2})zC(q��uf��J�ݘ�b���΁.k����J�6+G-�f�e�3y��1*����JD'���uFB�d:*@y����kP�5a���^�\�p:�]�o]�,��ɿH�o��6�#�\���S�6�X�.RS���d�w"1z,�V����k���h�1P� �\F�*k�w�ތ���NK���z�6FG���~,؂���QG;�Ӻ���T���@��Vw�@7����;�7��p�2v�=
���a��ۚ:��������ف�X���e0>���^�da,����u�9���� 7;k���J�x���t�,���sC�M�݃�s�z��ix�Q%rV�&uɹ�r+~�mì/̗<
Qހ�4����r��o� (�H�R�?��񣖆�F�jj��U8C��G�Mq��O��e	�M���G�|�/YL��ŀ�2�)]L�<��2��N�梓x�P����T�B
t%�3s�H��������7b���>p.����*�6�otLcYr�DR���~TT4���2dI->�@w]r�`��n�(Z�斖@�V���RKU�pwI��ӤqBB��ȞF����,<���u=���;K/&��F���~��.ߝ�ؤ���R�*L���8��nd�]���q�1��Τo3L:ۆ�cH9[�ܝ�ױ��"M��:��a�y��<�)yf�������
���3��⏓y����t5>m�6O��� �L�ݧ� `�_�K<Me�#��d��d{��"�����M�w�f����0�����M&*�K~$�[�VdPi�/�c�@�_dh� �2s�u$w�]�w
[g  �:i)���Q9bLGÔ�o��D��9�q��� k8n�x/j(��Gw�:���A���ۋ�,�\]�c�mD�t��o,lP���Tw��0��6���dצr]=]��5S����$Ui�n�w�P���_��H�SO��x���7�%�K�0�V�^�����׫V=_��ę��7�ތd��~%�����"��{|jq�Wl�����ĶA�#]�4�	���(��61M��'O������8�ba1>� ĺ�*t"��Y%A�4|C;�c6�t�����M0��]�!|��v�-xP!0G�eX�i�g�?q���i
}�Li������̪8O�e��A��X��g���Ǟ��F)lݪ����q2�^��l�)06j��r�J�y�s�o`T�1�׳��JSG� ��b��bv>�ϟ&�p5[o`a��L�JF�.l82!3q7J�),��*�}\����y�hzv�0�"!}��Ҡz8����ݷ�p,�KȜ &#c����&\H���0Nr0w���"=�VVw�8i�b@
�m�݉Y�q��X�m*��O�5��VW�o4�F�e��r �+���$=�����
��3��έ���ȥ�Nk9aSSS,3��	��f�Ns�86����Ү�����1�U=���'��rUC����BG{ߙwӓ��s�:�!���%��[�-W��2ʰleUUfUuu�/�@�����! u���܋��L� ���j�Z�P�`�Jy�����ׯ_'U�$�=x��^ۄ�ȟ��.��k��ڙ�;�;5�_JQ�ͳ�4%9��]ۗ����� ,Iwuuu�����(iP}�����"��p�s��eJɞ`$��
�d�bU�3����35��v-�ٲeKe�OY�]�么"���[����j/
��B��5��o"	}YM��A6�rK)BS�P�+s^Փ��S�E(�|��
gy/��g,`��o�1	;�/�a��O[#u:��D��<r{�;�^m+;��?�Ճ����/%�u���о�{G����(�eUT�l�ښq7�j�q�^В���8� ��j0�
�a�0�6�K2q�q8K�����K��)��>(HN�%A��v��)^b�B�[M��,TUPPؙw7�ϯ��cV�iu���4�>�~}�%�D����� ���f�{���>��'�0�:��)�:�25��G��w�.a7�}C(u'w��E�z� �,�z����e���|��G�)/Zt��0��X�>ۆ���W!5�
�$��l�?D�}�M�z��B����T��I���8�'*C�����z�Yb 
u���"c5����s��ˮ5޶\�ޙ�����jqpq��O���G|v��mk�LP�f� s�U �P���;d�0��ka� ��]0���?!?�[p/�ӧ0ȸz���aH(>��m���Ͽ�� �^��0��Uc69���	AE"|16o�Y���d��h���R�^����W] .Q�В�-� _��qP'�E׳(�nI�꧌��e�̲�D��@�B�f) *�b�����������O)�12��󇰨�d��2���T\-�J32��̙�cL8V��q���"C��F�*	����7��t��tC�tVf��M�|�"G�377w�-�G��5����� 8�E8݈(A���x�4i��vڡ��}#7G����Y6�����N`>r�ǎ��\��S�	v���~8���w�(ۅWm,_�N���
h �q�4�/��F���t/�3	e~����[!3"Qҡ�v$U?�i�ֹ���716��:�$�A>R��SC����Ū�5����W�ԙ-}T���o���|�����z[6#dk��O5���"����H��������sĤw�E��oC���I�;|�5̷��ѧ�ڳ��M��k��yI ����T@y���K�c3}}}��U�䩅�<�ga���Ls���Qg;+++��r��8_��pX�~=u�л�D��C�XX�w9bd����.A��F�ڰg����`�sc-Θ_--�6�:�e���^;������r,��>��y�����VB��y�LC}���x�eGG��1&��Rv��i�7���x��;����?�,�W*�FG�Y���l��y�
�1��;>�8zX�)��$�{7�L!%O�J�s�ςjbz��{	ƫ��)��d�oI;���,���N�5��BAp����\�+�:��:VB���D�,i߭�3�ԑ�gϞ]�:�Va�Sz�1$v�"_&B�kXs��I�|��h��=�`�Z�o(�VGO�z�q	�OKZ������o�������:9��,�%z�;���ob��3� �Cǲ]x�"��d�Zd���}(xE���:��ͣ��;J@�}�$S1����9s]z�z:3��A�7]i��Y�3;̉5I�X���tP���#�Ģ�I�MzP����W��R��AR�333����L��������x$�*�� ��^�Պ)�O�w��Y�����`!����^ŧA�姡��F~�+���M� �����?�c���CJ�W��h9@�7����������d�c��@x'���~��u@�E�M���ɫ�_Q�-��Um�4�!�Z����\�^���؍�r�@"���ȃE����[X���%2�z0��-�}d�8f㎸\ޠ�~�a�)Z�(��,|��07B�0��X�_��1�
`ǟ�J���;A�<M�>���;���=�+u�/l*��l���	۲B�<�������S_��	|���^?66vU�� dD~����Uw:H�w�?��b$7�4�[`t|�͝P���U�7o6�`l���=@�7��*�~#'�lG �Ӏ��VO^A�3��>$A��L v�sF���YFՐ;�O�ܡS�����ɨQ�üN����Q!�y����kZI���	�i��.�/�0�ȋֹy��8\�UQq�I9�:��:�
�b3C^�#�=v��E���mca�R���m�9���[��*����c��K��JKK31�g�������t͑g��H�> uX���<h)�ؐ��d�z��aB��7{7��M��A>C�xz���f���Qбj��hx�<�W�_dh��?Y�}R6��6�{ hh�W��, q[�㗜5�To�z�� t� ��M�	��Ѧt ����3�:RpP�����}=>L��N�- �{QR�9*K�����3J1���0VOޅbD{U76�8p`2v��B�7�N��?}��2u�:4�����ZvVm��V��oA6h�w<��uv�%�N�<ٶ�T��K^Nt�q����,%�+Թ�U��3�$W�%0����!{�@]�f J�R0v��*///'Ї��8���F���6$�=0:�+\ɞ��ѐg���A>��	7W�JK��h����	����L7X��3�L�g;�O7����q@+���wyV�ú�t��@,)>�������H�򧢼��uK���`a�ϧ?��D?؜�ρ]@̛�v������c!��Y�3�<�\f��.� ��o�# Cμ��dx�����㉊��U�j7�pQ3]�\� d��u��"�XvTvȹO��H�$a��!���ܺ�7��eCrT�"cc�5Z�*�"�$F7.����ʠI��,0i:�6"��������r��B���S �::�i5/Շ���6����(�D�T�U������ZdǇqCCC��	��_��?�w�)�{�Z�J~hʁV����6z۶kjhL?LuC�PZ��`�L���)�DUP���!# ��h�>��V�wf�`@󥺄�����:�a�\s)q��dBF~����X�R=LDpx�����L�����6���o�ԑ1o�Q���6��6��S|3�B�j�?(U��1���|�#G޽���DCf�mY�o1?T��4�Y�r���g��� ��Y
�����8h�����Ti�I�x�u�!�&�e�����.�V��a)}of�8 �΄�*'	ŗƌ�s�C�iK�J����r��!g�g����,~�Niu$�r�u٫���c��-� �y##CL����i}�DYHd2��v�� �^ja���9���\ZQ�Lڷ�i;4�<F�Г �q9�����0~�e�gj���A}.�ǙZ��V��ToW��� �O&߯�~׼�1����v-%?�tN�Bۉr��f����D;#L�(�#uO�K�'��i�6��)�K��<�8�cf�;2���-̱4�1�+HQ���n`�9�Ȅ)�oZ�} 7*�qG�s(��7��&)������GR$�����������O���>���w��r���6��i���u���JB��ώ$d��ǀ�����Ԁ����PRn�In?)*�E��	��p���=�x�5	�Av� ��/h]���c(U|X�aw�r�4�O�,+q�&�wy�S�s`N�&���e� �ƺΑJz2�y)L2)[��n�6@���*kj�O�4in��=Bv�-$���F	��� Y�8��Z4�n�m@5�̡�H+���	�ԓ����n�L�t��[�i)��e�ھ{�޳�����h��t�Q=�EG��U(�ZXx�5pT�-�����m۶堺�Y�<�u�݉5��!�Є+��O��A�E�]�'����X�x�aH����^ۏ�k�;5�jd�1r��w�Z�MO@CZȚ���P<љ�y���+��h�V��. �%�[�I�5�DQC�ײd��&���z�A#�	�K.�#���3Ϟ<y�vp�;I�R�q��,����D�[�y�:it�՞d�c�b�uf߃��(�򤚢��n�Tt�#u����b�����%r�
w_X���w�2r�F�ҫ8��5Eb����ڲ!3#������70�ؘ��{I�*h��Uy�ŸzrL1���yTsȣn��>��ֽ�Ej"^���p����vD�K��a�\gcB����YWt$�ğ2���gd�l<�,��jg>�?`$u�V��c��ܒ�V���,����9S����f����h`�`��Q���ͩ��)��<0�܂�Ў�=ʱ�Y�usW�^M�+]ۊpF6�nM:�ҍI&�Y�Y-���к���u�%�Gl� v?ǎ��-}�������D�mп�������)�$�g��>k�=M�ํm���dD�Ni{,���.�;@����x ��%�u� L��
��|>a���%���@=�Gy0���ݢ��]�ϸ�)������	4��!�-��8�ˌ	M�3<�Sr$�{�,YX�j�|�Jo���(��Ͽ��4JH�|���E]�<��8;�Kt'����e�WѯH�;;��$���|(Z �8���H���r���{,G��2D��tu�v�r��e��,u��� ��0ژ*��Sv�Pt���l�2sKصI�&�;��n����$ Ey�;3��|	J�1d�����&�o�]��(t��TQ/FO�n��f���_�
�ԙq�>r�l*3��B=�Dia�|{J�$�����Pj�BKآJX����=�J�}��CY�=�Z�ZE���3��뙙q��^Z'�<�ɚ����vm&W>��	�<ˡR�Pȿ�*����ɕt���݌���a�XǌIn�W+B������ఈ7|<��4R$�I����of� N�B��vV�B;*���&w�4��uf� ̿M����RR��0����u��=h-�C��C Æ�'K�T�BB��&�j"Nn�=�N�L���T������mu�֠q`�8k ��-���)�q���8mI��`f��r�г��������u^��[L/������F��RFF�u����9T<Wj����"D�>Y�d;�����S�2�y�S��KF�
�Hw$c�b*��Nh��2�r;��gz֡�ȃ��>ة���g[�h���@B�")�0MC�����zw+`���B�!ؐ�'%O��g�#ϑ���@'�s~�k�F�`,?O�l(`'��_�R���r��ݷ�E?Q/'}*M#��慰Z��{r�q�w��^��9�c��R0}��4 o�P�:Z$�y�1a -��1����+v@RdP����xĩ�,#�C���w?��82�w	�����n�d�|�����T��S�d$EB����y�f\�+��|a�^{��Q
'�{Ӭa�jZ8b�c���3{7$�]B� �Z��]/37��d�23�gg���1��sR�@t��T�5D;�u�dNJ�ϻ^5+����u�y���.,�L�"[� ��B�<Cܨ̾�Y]�<-D\6ɼzXX��km#:�ƍ���vn�>r/~ރ�Sd��Zm�x?�s�l3���d(�6(�Q:p,ی���e�/,!��l"ET�&���϶�
{�J1d8�oñ�d�\�9Z���q����$ _ħ��w��}�����U��"���W@�Ői�0L��!�Ts�t�^���PCN��ɑ�E��A^^ֽ{�W#�Tj�Ni�����-�Gӫ: �H*,�\,
�tm|Lʭ�����H�WF�A�n|C�l �	<sn�ؘ&�d(B�K��؝��fLu�K�f!BAkԩрtD��<�����f�+���r��nZ^��R�@�n�NLYN����ت�����>��h\X�����E\���?B�JI:/P����>%�K��9��ƪ&G跼�ϴ���.���g��7��n߼J�F��ʯ�j�?���U�%��/���~o�����ħm���V��vm����k���S��Ǎ�iI��S�n�3��������} ���/Z�(�ǧM~�+��B�/YQ[ŌQm��0��r�|���Eb酐����D��4|<:{�A���62O�N��n�rwj�\�cj�+>�KKP���;�y-G�'6�z�i�D!Z��X���=���K4R�A`|��GJ�OL��:khh�U���y)��H��ce���d 5��_��@�rI��� �Ϛ�t���D��O�}����&�.�I<� B���~�H�~wn?#����������bb�ҫպ�ۑ��a�(��z�� {���5��Y /���Gs�� ��!�ai�W����w�UD+�_?ņ_Q1N���"/�MV�x4����s8�v�A����2c���rs���3�Ô��wa%s���N� ~f1_;��������)�C���b7]xE�'�S�-����M?�Iou|���[��W����]r!P&�4��$-��n\�(�����~~�߭��jL>����k��j�Sz"���X�u�4���	ݯ ����W�:/@i4��d�PB��ĉ,S�6������r���s� Ȭ ,j�i*%���d���6?S}�i3/�Y�+�\�3H�<���c�^i��V�imZ�#��	y;���t|��c���,$���uw�H��;��s�u#�K��ў�h7}�W�wHZ�6����Z�(|`M	�<h�豈�F�>%;�^��/�?a�o�9�wEj� �&n�,��~�h���q��u᧟��s�U}m�R�V�-���H�0�{�u& g�nbjz��3����d����s�a����:��X����R��/���w���v80���9�)�Ȩe?nf�����H+��X�bV�l��$W��I��Ͻ��pY��=Ym���!�.�0j\�'��f�������p٪��U�5���^=gq������T�ﾁ�����+5&�R(���0�*T���@TΘ�p[�	�=G�/�8?��j���~�=͊>�kw]��M�u�L չ50gw�4�8���C�e��j��i�̘�ͳ��y#��,�ԇ�`>W�q�9q�R_���>ρ9u03��7���wã̘���VR�>��WYW�ԕ��CG��BS��B'Z�� A\�������Qv���T�%�*i�eu	j1�b�F�Pq�@A���(� ��u�	�>p��}��ܳ|�;��{�O�X�P?��t�I�a{�Q�~?c���;�ˊ)��ɍćtV;�.��f����^���:K�t�����B����~d~ӷ8WB����ΡdH`�]����P�+C���qYwMdz@djw|0��6t�իW��c��0���R��G��FP���oM��mf �EY��$�Ō�Kc��Ż���9���ݓ�b�?|�Q
�_��V�:PRb�pH�ڧ4���2G�}*��2����g�������V�4�[ ����T"�n��F�C�36C��� ����ս��k"��-L 3H@8�/�s'S�X�]�"!���_�	Y`�_MW�,���\<�F��cnl!��ʣ;k�GD!��s'�ȑ#.�`���� ��R�=^�`l��~��P=�}߄J4v�\��y�b�Z4��D��0`��o�gI���;gŻעmR�F�;��N����JJ��ΎY!�e8I��è�ą���w��G9�V��_�ݶ���Ũ+��]�e)v������V!�=�n(<�R�#��h}��Դ��䌞�wI���$;���L�:d�<i#Sa,VnaϺm�H��=�a��T{}#�(r~��oo�| ���0;�����k�M%H:R ����GB3��Z����8��Q[�X�W�mh��%1Ke���q����;�.<y�u+ڐ���o����=x�4����.�p)�R�xW�����C6p���uO>[�Z<k�c���#G?�o�o�D��;�*��c�I��_xR��sF"Y�v�4����{�>�! �-_i ���˪�B�4�R�5�M��k�e���Q6�.���0-G._~T4v~�W!���m	R:�)�r�n���������CXMҏ2O����G�pj��V�Z��b�]��`4-����?b��]���Dtj�P�<2]��U�-���;gb�Gr��(����W�n,B�bKr5&=�y6����I��#l]q����R��Z(���-z����	��� ��{��LUe�f`kB����O�)S�*�x?���R�NEW)���^�♼N���ܯN�v�Z���S�f��.b� �j�Z�܏��<�%���r��`ΰh��yUأ��eꖑ\( �u�]q�E�@�h�kj�9��41K>	�n���Ӎ�ƣ,)[�����^�_s�j��`'"@�Wmp�]��b�
(X6z�����՞]?�A�0S�`$|���Vnܛ��8$�I�S����\]�O:1���!�C�7U��/w�+	δX ��Kt��ء
��J}$��!���B��k�bF��q1�UEEE�h 3iN����JM�Ʌ/�2l0��r���FVW�k��L���Qq��l�n<�qCG �7ۡ��?-..��r�g^�u�Ɣ|:O��HP,^����~���P�>Z˛~��JQ(6��4����>�?���zo1��O[���t���$	V̉��e�a��i:�U�� RX��J���ܻ����5�*����pLB)D3k�i��ZV�ד�COq݄nU�Q��Z�x��m�i�,�Aޑl��.��[/�r+�j�|����p-k�y� "Bݑ�a``��V7�E�;(�<|����
�jl�@N �u�Z��@�u���`��s@�by�y@Kl�b��OԿ�ܶ��r��l��'�(+��O��GM�%���9���-j1����0�������Q��2{���Y��n���3� ��Q��.����yyZmc�tҫ��wbO-�A��"�kӚ
�9�+���&�����}��a}�@����4�zTep�fT�<��ď�w�ܳiS#�9lQ�p�|3�*��#7!�n���0�s4�4Å���y�T���qu!hߔ��Lk�}���ǅ�^UՙS(���^���|�x7��U��Wr��|A��(�B������ၞSvEy�ט��S�?���ux�!�-��GW�^$A<�&�Xxy��XKol�A��T��!rFh�y�k�:N���o.�@��1E�����Y0R��H52e��S� Ъ��xҟc�qM4���-L=�%AM^<d������������l�T�hg�i��'�H�	^j�{&�^@/do�܀ :�t�Pg��2 �6#�%�+�Z�s?gDa�����y~�F}���OA���� ~�ԠǷ��J�ہ��]8��k�������u�����+�1�Y��d�����'N�]�]�7։��!������G&L.��!ЬA�b7�s�^/�x��Q�,��"�pߛ8C,�e3����>��kf��FcT�ݾQ��Zz3j��b�z��jv�J�z�)��W%P/Z�*i�iq�
N I�C��k�����7
BS�R	Pc�j�ׅ��""��8e-0�� ���)� ���)�u��eHr�g	ԣ��z{>s��t��\���H�	O`��xbe[֘��x�k��N�x����*v-뽠��n$B4�=�[|��va����y�S7b�V�&98b��%��ɏԻAU�k��m����<�p�A��}&�L�8�[ox�>'���T�]�����V���Mn;R��q�����`(!,է�B7��i�h6d.���/���ؙ\�������*k�0�߄�Q����_�
���)��Ho������Z1���Pp}8�W�ye��Oڄ�2�t�@�Bڧ�rYf�ծ��a�G��B?�8���ě�eL����?��F��#A=�m�	�B"���)�"��=�,B;NXd0���S�m�GO�K�����,o�`Z��s�w��8ԖG￨�y�5R�&Hx�-ۮH559���>����xJ��e�Uea��+�Yꢏ��-�q��������w���=�Y	L�,Њ�4�wG�n�Κ��\5KJJ�I�!d�3�� ��0�{����< %�UC��ȫj$]5�L4h��:K�'��sR!���\�@��ڙ �
�����'v�d���:ko��a5/ca����!I��X6d ��Ȟ)ɼˋ������
Y=�44����/�d��u=����v$����.�j%*�f��%��1g���Bt!��!�UOzw�Z�V^��y���'�v+-t�W�9�[�qԞ�H��~>Ϻ|��KAJ�${}K�cW$?
vt7��a��t<J◑�����Ҕ�2�=�����iҸ���~u����&8�*���yT���N�D*ډ��L���;�F��	|5}�c�!�b�8���&CL���	o�~Pc߯*��/��`�PGn@��I-�ɂr�m�]Qs3R/�n�� ��qM�k>��ء�e���%I/�L�O��iX_[�GkP������K3��Ł�Z7A'nW�Go�ɼq�ShvuԠ���Ҳ�>͏
��e������Sw��� ��|����C*l{�I�FvN[���h<�2'�Qn��-���u-P�c�����]=4�	��T�'<X�Q5a�R��D,@D��t������=_pI6�����l�"q�t�g.(Y������$e���x���p� Z�ftҲ�k{�g(��}��U��gzk֭.�kۢX�0�5}���bh-���݅�����jz�^��|/�vز�|�o���Ƒ������ PK   6��X�G�#  �#  /   images/e0d0e70e-96b7-4f7c-9039-c9e958c885ca.png�#]܉PNG

   IHDR   d   E   �C�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  #/IDATx��}y�\gu��U�ګk�]�j��VKVk�,�H�3�cb���g�1�!!a�Ü2�rL �30��ld9��&��Z,�[���^��Zյ׫�����ڻ[����\�������{��}-c�$��L�f�#� ����R)N|����_�KH�#~��b)'�:���}J��!�$cnW�`�M|U����b����;���w.�9�����{��'�K�o.I y��B��,e%Vlm�`<�D�x~��'b�ȆP4��D�h&n�t�s ,�ݱ����8����4�L4%�5�*!K�y]	j��+X[n��]A�9�k��q?IұH��w,M *��,��1q��LG���y��ٰ���ӂk\8I���ͥ�P�l6�F��p`4��Zj�&:��o�ֺ���#���)�G��WN(*:�t�C\m�C��?�9:�"z{\&���;����F(i�D�|qII�i���߉�C ���[�o9C=��{97�e��8d�Ű��u��"1s#7�Ў��B'}�Lp�{N�� ��"�W�ѥ%��)��Vz]�w,����?I�F�!����k&�g� �lK;.�J��FD�,E(���C�E��&�yۯ�G�7����l:���8xb�s�3h�u����Sx�]f�M��z2Y�ɬq����#���g-�1\6KP��~&�`�YH�F�^�zs5C|?���v���`X�
�$SU匢ĚD�+��)&���&�rR|ŧ�8�q;�u'ҙqj<��ۛ<�S'S5�L�%*�Ni�gzHh�7XzG��e[9~~d��\Z�y���EI�Ud��{��?k��2:�����t���Io!'��w.�IË}�H�f�ݘ�9fi?G��&:�ь9d�ms5(+��s���ӎ��s����"qS�p�Sd����t��d�Ք�K����}l�4:?@��LǨ(�X8�����e7M��	IW�$�y�;�wp��o��L���w�gi&S��B�5����$i��ZWL �{Ѿ���<ݹ�c�j�62W�M�j��01��,�cш2�.6k&��*#c�1AQ5q�OO"I�@@%	9,��0���/D(���0_�ɺ��ff�x�k���:Xh�Y��b6�	�/q�}�6���?����w5`m�g���'��I$~?�?�:�:;�]�����:Tj�@TGm�c�$�0g�8��΍M��D���#c�Pp$i�����������Xԕn�C�V@L�F?#�"��ĕ�d_��?X��"~�u�>$>tM����B~��k��ٕ�ޘ�~����4�0�)�jD�ėn����h=����)	�^���8����zo��Á��y�����[-p�^����M��5����������A�?uc�^KҊ����#f5�`�d��ؽ�/4�n1�#3l3���?Φ�f��Snk�Tk���3�y%���)�iQP�
��҂�r�p7b��w�ۅX��H^B*�Z�ndY�a��H�g ������9�K��WK�k��:�0Q�[]����5�C.E1w�Ş���kSu��@�n��d��@$�&jDvd:}�����ϓ�c����29G+����gM���`&M�wY<��c����-�.Xe�@��]�YGJ�/<��x�Q����L+#�L� ���԰�&����]�v����M�����J0���dxF�nq,ӹ�
��u�]��܁Ɉ	��Cm3В6tLV����lNz|�Ԙ���&b��	?�]c3�Ϸ�G�=^=������Ү^ ܣmr!��4B<�tp�I��ts�D]����O�U��(x����R�×�q���������L��.�r�����{�z�k	F
��,B�<�xDz�$�#d��l������*&>���q�u�����!+���u!<���tB��Jp"z}3�)�T*%8Cf3E֖+���S�_O%*�R��V�-w�S=q)����v�W���lQ��߻�; �H[��\Uwe5�[�����/�����8p[���I;���|�}�x`�{(@�	�D�n�����K�
ĈRM&��2;����&R�S�d�:�I�5�:(����Ӂ��@8�yH�5,LҒ2�"��,6�Z��aC@�wc'�j��	���������$RC|+qq������a���l���8K���f��U��lq�d& ��83�^M�7hÔ����D
�!)�:����	�d܏>Sz�t
_7��QoE�H���R��FJl:��w���dEq���F�Qy0�Y��'bBRh�NQ[��LZϖX��}��������C�� ��=������uT�ѳ^����T-J���\j��ĸ0e���hhlµ�n/47�LZ��W������ݤ���d�7�B���u���O�L���oȌX�UR��^2˕��aZ-!c� �x6;��o�u���xq(���1TN<Hb$����?���L�����S��a/' �'��.W�(��ص�s�V���ÌN����<���22a�������~,�֌�{m �_��?���A�-��� ���;�ɱ��YɧX���q	������O�C�&j���pc\4��%������t
��uB4\�dn3�������a��t�|�(J�m��4��W��^L��ٸI��H�ش���D\��i�o�i�&�m�_֕����O\��ۀ�C��uT��3K���R�_�9���[��.C\Ѳ�3>A_�D4��� ۦ�"'�H$r=�����m���B>F%mS�vF2`��6�tM+���--غek��4\���I�4�N�9i4+5��]�1s��Za���5�5u����N���??Y��h	�XI���ݸ:�Gqs����}3�z�K�Lԁo�܉�����b7y�+- ��G������P�AH��t��
l62X��
�+܋{w����ʟ��9�� �Ɉ*�����8��q?q[Z[��d�и�h�e^\���c��J�D{ka��^GUX��kP���o{�f�Y������DR2m�4���g$�,��"gS���ԅ�:#"�٤�&dz�,���\�%EZ400�ᑑ?�"��D*��F2��/��|��t
��!֐�D���ل+�������w�<����m�C�b@*]��Z�j�%�'[:�����n�G�6�����@�K�M�*F�RE�I�Ø���B��d4!�H���c֘$�644���F!H�Q�PHP��<<���!�~jHÜ��ڒ	-��,�贶(��=�cK�-���1��1��Y>6Օ�c $�{"	�؁?��]�M��IP�}~d��	��Jj졞`������.)`�p��'O��^cڑq��X-V:�
��)]�-�8�c�ee���a��m�.�֒v������A��h�(�_�rK�CR��ɺ��ma�"~�C=xc`�{~פj�;Fьt	��ܶ���]G�g���i?��Bߠ��)פ"��@�9�R�6Y2��Ss�,����;
sO� �+����ҍ1x�#��n���R��D��8�`/u��N�D���B^�ϫtF�Z�$o�3Y뜟,CR�;3�L�`:��NjB��K0yS���	�~���ӗC%2����@X�C	+z�>X"25���ct��/�a�wy�.O$p�-Hf06�������b�K�x��(ư���������Q��˾'�����>$�`o�&�����8�7zI�e<I�� �'��O0���������&�Q�]�P��D���*��6G��\9��c��j;�k*�'�ݙ�)0�^���-FH���6�!� 9��o��*�Tf}�_6W��1�� ��t\�/���%qf��N�H�,�咾z�^_�׬s�Lf4iF�Ӂ��
�����&\��:��L$��Ѩ��4h�����y�r��tL�o��f�^��|&OJ���za���-<X�Ρ��*
DE��
�ѿ���o����p�-�b�"�֊q���wr�-�4'q�~���f��Ћ;�Ȝ��֩�0���r�0��:dS��/����]`�������k�g�j��B,�=5AyEiIV���EE�ef4��D*D#i٨{!��S(&� u2׈%����n�D �`$�@�-�ϰ�~����G�NO��ծ�g?�I�ҁ��Ut���=8�ܿ����ye 6��<�%���dsP+M��<041GF��H�_�zs�sR�^qbq�����8�_h�2b/����"��/�`Ok)�xu�րWΎ��F��?$�;I����޾�S�{9�=8:��	��%8Ge�L"� D��*T���[B?����9A�QK['�n#�U{}Z�o�%"�� u�`�J��86R-rZ�o��ﶊ���ø�ɋ����c���B_&ػ����K�~9���ר���F�N�����|&��̧b�\-��Z��:nl����L�,2S1񟷝�z&!gN��3cM�^>oW���Q�G�rF����D��%��W���IE��4�+��
��Z�7�����1�/:�QU�����iIaMI��]����ee�t����@��
����P=���W1�'q�R/w*������K���9KCM�¬.D��ѡtM�j	JU��K�TVG��*���4ޓ�l6�ϣ
���!����rĂ�b'q�9Ur��)?q\��������11>�#�Ym"����6��yYY)\.�
�{cw�;@`��!48bxűQŌ �����*")X��,��p�M��5>G�y���/�X��"2<�O�X����]NэMd1X�_�H�_�u����$E21ip"�������T��4|��#hjlĽ��Q6c̹��-�Ez��F�|�F-5ؖ�1���6��C��ݗU�-�r xwC>�<%
`�8+���%=�"؛�v ��\h���U�|r�9v�C�Q���6K)͵�&KAM�dIq�#Q��������6���҃5���&���D�=?�~�l!����ܘ:;]�"P ���LN������Ѥ3/�E����`]�S��N�$��2��bs.���`�ҩ/:��Wɱ���Z:�����U�e�������sY���2� ó�2���,)HP�908(L\�|�h
�}� ��4T%�X$$���{��H��/2YwT�e�'�����x�ח-��R� kF�ߎ��Dq��r:5����(R'�;'��YS^
�U�5���Wɚ�W10�D�%KI����Ke=�L���ٳ8u�m�]0t��5d�����ޒN���^l�ؒ���d�^��&�C�J���Z27��z3#A2Y�xC���&l%�\�.�eS�R�:���;pq��(u[((tc2�D��FJ�n��B����w��O�O����.K �Z^E������Vb}y�g��\�9M���EIII�9}^YQ�]�v�n���@,"k)*nȌ*�Xa�_��aƭ�ޓ.Ñ���#�ƾ���{6\���=uI1�B�b�ֲI��f{�!��
�!q��L'.��.p�[Mx���j��J��|3��mo�z/�9�]O&n�(�&��w ;�0À�y��\�����������Ŋ��\#��TWWQ�Fl_�(C��m�o��~I��F�a�5��#oޔ{�� �[Ǣ
��d�|������!v��"��Z;4�{0��B��.�a&�Z�C��t�H�`��ඍ������nh�!Y�	������}q������V#�hʯ4�Oܸ�$���n��{3���t��C-���c���|UW�b*ҰwkHkǢN�捙sK#�U���757���٨�V'u5'�DR�\��V�����v��:�e��н�l/���^��2�K.�v��(��:��̩t�]� fP���t
��qN�8�#��m���V[DkX��J��U�h�ڵ�XS�v���!.z�� ���(-�!��񸺚'���$-I�x-�|��Џ�yfpn*_��̷������1&��J�S�Qۦ�n�e�<3�� ��5����n�����ʹ��%�����CO�.'~߈'~n�w�_j��zfP I�p�|���&�V�wc�����Z1_u72;�GO�EB���]F�a�nm���"#�]|����c���Z�7΍�E1��<�����i�jb�l"���W	�Zcy�[��/������D�tŦ*S��ʇ��mֺ�$u��6c��&�]S�#ߤaBj�����Os�fR�[^�H�U4Tʢ��Lwk���r�{����Sf^����x������wb��V��3�6���{�=���jˆ�:[��*x̃�RܐS�ӈEc�P�^r�;�Z���ۍxA2+v���쁗b��8|��C\��S�b�+C�k8LBQD�O$�f;W�O�ᦈ���FDT�6��_�&��Z-���<��׻��!��܋����j����v��P���ك_:|==���L��8T/8'c*o޷-Z��i"��́gEݮ��_&�.&H�W���Ϗ��{��\-���M'2E�b/x@!*<�	EG)�<�Woh��<eqz�Ybg����g�������]�>\gR�yK+������/��Űmq
$󝋩S��
�D����&��3Oʕ)���Ր);��f��{PF0<���=C6܌*�������6^*�̊e֌-�C���q��7�u%!����]:'#��<����u���o��(ט��LĨ��b
���킓"���
!�7T5'(�d���N!������_.i� ��(��3���7\�ýA��s fYF����3h�<v�4Yvŕ�K���t�H�_S5�O^{.�%�Slsݿ�]��6P|�H�+2�b�@�����sK��ϣy�n�5l++<w� z{���I7~~�0ߌ�o���h^��Цt�r��F���O])x��|)�,�oR5��N���3�"�̳2�+A���w�Z7���8⿳�����<?������������I��`�Ȣ��a;gR%.R%�DЛ775��l�dd�z�#��T�XG��]LN�"��y="�7�|�<�P$9FC�����z|�!��H��$�u��YN����3�E�f-�����n�Ə{�������)!�ۈ"Rm��u�����8ї��7��5!�d&5]		���e�7��>}4��+���m޺�`�(��������Ygo�c���X&p�:�Xt��&����w��.�����&�N����H�b 䞝V�Z�w(�4<�vīqv����X�<�S�"����`����^�I����q4�âLRS�8>p��B����W  R����0_�ܰ��~��z^�˔)&�3NQ2uG�Z�Ӯ�iS:>	��� ?�K�E\�e:��4���!�:Q���Q�x�VPq54���l��
4�,c� E'�F���[�Y7 %�Eg$�p���8-.�%��rI��?/�$�m�e�1�lJ�q#@m�F�P���y�w�Of�9�G1��� .Ԓ��k␒3��c�f�mcn�i5���ݖ�f��x=sS�$��A1���Ϙa�w�f�'� ����y��g��^�	����CkU�ע�̓8{����r�D��mx��?�@�9\���M��Ճ�d5����$���������\�p<%���s�jz�kVE �ULܳwT��5���ԫ�*��}i m���}�q��2'�C���Ћ�����c:�9�jW[�bذ�����&�+	�S'<5����QD#�[� ���^�xG��&g���Q�\V�
���>�7�P,%?�(7�o]�+O�5��@~��+�y���ֺ�bLB5�%6��{+\>�jS�@R7�ގM����[Ǆ�g�xf�u�~\�@���M��L`��b̚"��<����w/#op��1���yE�;u�d�P������e��V�Tޯ�L�����/�?��}�����N�`�6��p_B��J���@�-�s�����{�Q���<�C��N��x��L���^��7M�<sG:����K
k�}ȭ�ء���%M����87t�19���oS�Ym���y�%+��*��/��CDY���u�}`��W �l��`�aJ��t�[v1ET�b�5>k�����N=A�Q�� Xհ��#����̲@�1�-��$��"°�g8����(:�o�׊WGk���%�����ypa�ڕs��ٻ�׽2��=;Q�h��l��;�1=s-�+�D�녶�⊲�8��u|Y%g��Z9J�-������\&Q��S��Ge*E���ŰH��A*<W�=����r�\����5:�n���4�H��C�Z�!���v��裠�o:o)u��XkBk�\�̾e~��^hg�n�Ŗ�o�w.�pQI���sbe.��\8}
�w&qf|ɫ�]O̫q/�|�R/Ă����/��Y�ɽg�)��>C<��k�[��d��	��0z��j�D�o��0i�=�S��t����u�&���x�HL2��Ꭿ�!m1
���ԹG<I�)��m��`��o8Ϗ��u=2!�;�'����#p{s����5Xᱢk$�5naO����X��)��yȳ�W�N���&��9C�9�P45�]x�KsEu��
�e{�wmJ��Y�z�(k�u�`ďաK����x�_(�,X>�$:���?M�3v��wq�'ϒ�d�0j�ucd:.Fֶ5x�v����r�/��ܱ�9{W��
b�x��8媃A��X=����	�e��/F�������9�\?�24!��Y(���ָ��OK��	�����Y#d1>�-$����w'ys���`�r�jPI��z�����o���A�'�ي�6�Ό�qܻ���*Ь�A�� T��ۨ@��    IEND�B`�PK   6��X�N��C� ~� /   images/e23486d3-0dae-4ef6-ae24-86700798fe45.pngT�TU[�=|@Ri��AD�PҒ�tw���[$)	�CwK#�%!p��os������1{��Ĝ�Yk������/�_�@ �2* ���������l����U��A1~Fu��r��;���u[�~~I�"��������������feg�lb�`�f�d�v(HQ�>H�W�H?X��Uu�A>^�7'���$_FJ��������o�Ua���(�~$�4��'��.�rU���w��HF�Vn�3}�@0��������8��Q�0��t�C~x	����������X?�3v�f�F���u���j�z��Oz)�(?7�4�5���MD����Z����o�0b���������z��ԏ���ԏ/PF�>l��7�b�Q�r����i$���rTY䡧_��.֊�`t%ɏwJG��[+vӔ���e�1���)d9��jJ�<���LUܸ+����~�B`�Jl�OT�C���z�q����ݻeYR�
�DG���P�c��]����p+%Ѱ��)�@�W	�,g�ދ0� �A�o��+� ��dWH��.$���<]�z�����t�8�ų��1���p9���߹���~xyBn|�g�蓰����c݉n-���T�嚄�z#쿙g*~X�k��BW�A6a����=n��|dj�����>r�͌�7h$�I�d�)���YC��f�c� h7տ����������)�&溂��θ�>y_N}A��!�MA��A<�Ix�b��Ǻ┮�.Q���/�S��PFRE�&��-د�SfXl�?��&�3@*���&��K�fP��]Q]~~c�B,&��Z�����M�Ӏ<T�_B.��~�{�AfX��TBjV�O�B`%0^Q*tN���m<¡
����lK�(Җ�����#%�*I(�M��V�G�Ѿ���oy�������\n����t�x��cq�F�8��M@UL.)UK7����1��������
�J�� ��0�ý3d�gon��,��g�h<�;a���j �-|J�_�Y����3q�/BKS8g�Q����tH��oMɨ��E�;v6�j�T9R��U��l�z�3�66��V����H`1qXJ�Mx���
J���8��HW#Gl��,O>sLN����|0�x��ct��eq�]�8�Xn؂-��5ņ�_+���l1�ϣ���@8��*&j1�P#�ǽ�)�'�O8_a�ۣ�1;��rT�j`��r�xJn�&X��U�ac�;�0���UZ�q��������Cx�e*�e/����k]ұ�AWA������}t�`�E��0�l i���y���^��&�iF�=��J ���"��E���#%������ �QכY��V��2�pB���g����p"�]'K��'Z|������}���P���{g�t��I�r�i�
 �OxsY�25y�F&��UB�򰀚����/A-ދ����3��Тgm�}.���"�'�Gew3kכ�%1��hV8N����&���.�>���$��\�9�b4o����Y��©�,՛�Te�p Y�Q-�?xI%�d�PB���ԡ_���5+���b���%��.����tY�m}��w�>�܉;�2��l��xDKͽj�f�|Ӽ��˘̺�Y1���8�O��@�{����������6���\.~�&�~��T>I�I�l��s��
�����t���9Rߴ���G9.m�y7B�pr���Շ��`��fO:��4VFw�M����;�Ѯ1vcWc�Afy�%o�W��Yv^��ɪ?�,Ō"�%��|�P��4T0"��1Ȳ�A|�P���L�w�����J��~1Bu}g�3zz`����y�r]TM�}�	��|Q�j4}}�������\���C�����FQ�_��}�Y�W�㷮��A�RWh�^�Ks(tK��:�SK�n<��4y�%�3n��#?mP�G�Ȃ�BW`�0�v�/`;2�@iɵ�-��6>Ԭ
~d&8��>���H/�X^3#%6N��&����T��X7�qB��<$eI\T�-D+��r��5��^�e7�ݞ)�\��&4�~�����w�l�:�t˚�P~��[o�g7��pf�������	�������ˮ�ЎU�;$���Y�۵����RGʮ�eb!���]L���[���rsV7�h7%���'�j�3�f��?�&��� ��A���նo�M{H�+/s��m�@�����/G���Y%��py���/Yi�G<_�ztϧ�9J��N�P,����}oD���㓏G�"ľ\w ݵ�F�H�o�/����r��L�bR��8µ��aI���ɔB���44Y� 0�����@����u3寛�ڎ��f���E�"vmk�������Fs���w)\��˵$%b̜������<����k���39+	0�D��ť��Tu4�c��yt�����>��c��]�s̛D���]���9�vh��g)ìa��"���\A���B�*�,Ƈ�C�# kj0�)��S��IY�b�t-�=��Wr���Uu���0/#�hL��l�^���v�`2IT}���=.O���KI�S`%�N�fo{n��1I%/+���W	�Q��(�
4+�w��/s{((
]ÝS�K.�L�3]���CC�BJ䦝��5	�t~+�
���:~�Ya������E�GG����?u�d�}�ǌd�"��ʜ��C=����nz�����xQ��ٕ�5Л�<���2]����k9���<fhO{�&܆1�܀��}y	@������.��̩��M�[�*��e?��FF0I�&��D�"hb}plr�MHݺzy�++���k��p�I�F�lc4���	���+�,�T�/LL��2c����kʇJF��x�:���>��Nh�2������M���˿�7�(����eB�sci^��sR-�6'��ԄN������B2m�������ˆ�����_��ݭ�$"-��z��8J[&�������U��6y���{�UP���?jO�d����
��V/���s��^�u ��Q�p�T -N�à�oJ���YΏ��>)�����[���	^Ë#��殖�B�х��D5Î��o���<8g+;�_�>���=�i:+:�`���V9��<\��J�
�����ç�y�s��_�� ���%_v���Cۺ��{�>����F���V$P�F#+���ml����j'�6�"��iě��w���7C���?y��Dݗ�T8�4�� R�oq[�ߕw���,u�L/�l�J�g�����t���Z��yo"o���i� �4�1�6�c�����l�^'����������s�����R�F�"��GnYr�b�t��|�ߢ�Mg��6(����f��y���XF����b���\��t�;�<"ҵ����"R����ȁ�����Y�����lF�����/���D�r|�v��M��^�m���_��������&ll���*�،�7�������x[����֗�w~�7F����4�6*,��P�ߺxg�2&�b��:@g�I�b-@�'�%��)����R\Mc#���[W��ӂ���d�M����nԥwM�bڍ�li<o�0��P�C�xl>�#���zLp���(p%bSJ)n�Ȑ��|����4+,������!���V�g��bCZ}B�@�t�9zw?�9��Y%��5Nۏ�~>�Y�?��=��,l�C�*U���d������e� �1�TR��;m<���&���Ze2�$
�*&���z�,�^oQ�X$���dL@5~?gr-������n5Z=�߾#|�3	�Q����~\H]��!������f�(�f_Ԕ@�n≮�Ͽt�U�ew��V�؏��o;t�n��D����*��%'�c��[6\,�^���l�Z�\<Le����m}�����}$Q	�ӷg�0n��Vݵb'���G�d�Ɔ���x؆o�#�1HP�>{L
Q�:"P֑a���l|�T��Uid7\%�Y��0P	՗���jq�&�G��{)L�$��Ԗ��j `J�)����ӊ*�oD'G[��z��w߆�`E����$��ʁ��a%�^��3w�V�H� �^H�N$���z�]~%�0�,
���b�FN[�Bj8�
rea�����֭��\0;r
�~]�- 4Ѵ�q�?�vE����_}kj\P�g���ʿe�IxǗ�D[A/(�6��3l�8�y[��j>-`!x,��<;�ϙq�q_ ��e��7��2���e�]εyP��x��{!���$�'$Ƹ���P��T�
9��=��J�l}&IW��#ߵ#�~+�D�b�2���>~%�����	;/�L������/�Xp�`�B�7eF���<�N�������{�a����{&�_O�&'�܏��W�>V�pp0�7��}�̓r�>^��\������]�VW��������(�ފ!CQ�ᱮ����P%(�X{�q�Q��/��Ҕ�05X��ۅyA�⽧|��DZ"��O$����~�_X�n�+��5|K���,���l[[�$��JH�a���詫���H�"xsl+)	=�a)b�i�2Mkd�׬�m|�K�D�A���d܍Mt`��Ȇ��pA�������3�FuＴQ_��=	/�̘��:��Ά�f��>�n�wҟ^~4.��]_/��)����Y���~��9�7&J1����z��w���ä����(�[͡�?��y7�����_��������<�O�U�*
�}����:�_��h|ȩ��s�OP��^��� E��o�0�}GϤ�~|��@���w�A���ÊLI�����wc�|1=�O�ܮGH��?�_�E�
����X7���x�����G>bL�]>��;%"���᫉�0��V�aY��D�co���I����v�12��[Xrv���I�l��� w3n�jJd�{�X_q�P_Ĕ���\�Hz?f���1I�����X�Mg�Y�����D�Ȟ��D�tV1@�G����~�j�\8������������g�z�?�rl�/���Ԁ�.{6������lY�x3e�2"�m���Y�{KL5^�Nk�#UV5R�X"~!p���T�W�wYU�Qا����zǦA?$�\�"�BZ�����P�f6���K����,z_���芄��u��4��do���uT	��Vܰ��u�9k�Q�W���E���ضiv/�NO��{��Z-��8�q������#_k��ܤ�����
$.�ֿ]�����YQ*�����dtT$h�~��{����<ť?�����h���_���|�}���t�k,�D��
Pu��S��,���OA�?�}^ R�mfڤV������g2�J�� ���E-R7KN�4;/_3�	{u)T(��e��SD7��,wR��P�0^ٔQX�;��y�\'n��6m��jpUEp{XEi�)��B]sT��=G�������+(�4�m�'�4�*p��5��R�+�^�����
� /,U�׷5X�N���*���]�Av�jn�×�2��4�iG������6� ����8��$M��h�?� �8����> ������dG��V��������Ä8�'���f���O&i���ʩ�����;��1|�t��}lg̀�yG���e�Y_ܟ��x�A&4�a���� ijJ�N��TM��¸[���kOU�k��.�����t☐se=�Ev#DX��O�b�u�@��ԝ�:��gaJ��s�qMP�#��ؼX�~��F�a�3?۠T(�/ή�4�
�#s�_��;���Ā�L/X�G�C4*",�՞�# ���ܷc��ّ��s!���FŖ���JX��8!a}DK��g��ʡ�P��V!�R@���7ќ����Z�.��+���b�+�E*�wC(17�8�*)Ľ�8���G�vRP���:���r��/��9Xik�W1>�WA���=�%>��.��o^��Ǯ;�oG�[����U�_��ΎRszM/�B�d<��S��"];-{F�<Q�����F.>ov\�yCH��k����*f��{�$�ZL�ukJHl�Ե��nHlf�|n�|���M}�0�b�x�(^���v���-�|����S}�t�M7D:��;Ŝ�+��QN[��Ap{zW�*�F���z�����	wa�uzM4�W�. ���%��`��@�}b9�p��D_��o�
.�8��`�1�������:��i�?_ݏ?�@���hk�Y�V�-���>X+�������A�~��(߀;/n҄-:y��a
>�>�\޿��hV���܊Q��Y5f+~���嶯�r�����r(p��^�A����)4ɛ���pBoݵ�F罓�&�\�?��ʊ�뉢���ugD�+���k�㾍�Ȟ2�i��S�]&�_�i�� h�T��i���	�}艿���S�,��:�Lͯ�}ܗSd����R]2	H���X��IE��ߠ��<q�`	:k��������Q��}�J�fx���s�l����6hn�0g^'����2����+�>}	��_����C|��p��
X�w�X�-#�F~���!8BF�����.>��|��o@St�q��/����m�5���S�]/�~▰ve`�2A�E%4n���ؔ9 K�}lċ�qC:m� �4�e�~0�өU��z;��`^���޷�N��j���h�{xN\�����n�pVeq�\�-6�lNZ |#�XÕ��� ��'��qϽ-�y{#���m�$���o����r���mq;����߁&�i_�5���g���t��w���"��h��0�Hߗ��/ڎ��x/)'9�� :P�/�+
(��k+/��u!�'�^%g�����Z��3��?���?�/Z5�Y�!��
+�Ϳ���4k.���&�U]n���=�����?N�g���s��y��z�������wb�խ�'�g7y4.?m�>�xD��CP�/�����Y$�t]�5R6&�t��F(Yo�p�����9N�־f�k	��Dik���j㪀�V��E��.ɡ��MP�#)s�+�t��ޛۦ�vq[\+r��!�4���H�����z��&�W�)��cVk�]��p(�(|Z�ڕՅ��Ύ��\'���#I:#ŋ����ٱ��[��dPT��5��w���e�M��P3�������K�l��ޮ9&@oܓylD�\���9�^^�c���^�I,R��r�A\����L�l�K�6����*�O|�b:FJ8C`W����:9ݭ���T���Њ��R=�/6�i��l�}�	$��������iC�4�W!3��3c�����m$����o��Wx��ϓ�.ꅑ�"���Ȇ(k�^�h���:����ͳ�O/��ج��IE�%'=͠�ݟ��7�sD�o�%���^��j؇�.������-��(�`G�d�D�L�����j~�U�V�ˏܱJj�c@ut�~@9�N^r�Y'��08'}�e�g�rڗi��;Ů֒��W���v�̪9�9"2�6�p'�[�Mq)�P7a�I�t[5���>�a�+��J[YRR��z�xDG�m۵��yJ�IG�a�
��=�b��g��B�S�EH��+�5>�(׾�أ͑��9 q�U�	��]~��#)��Ȗb+��?�:��i�*��C;^ca��ļ`�IF� '�&��\���nՅ�����������e�@��̸d��������x<b?|�˭�c�l['�1�94-���5�B��ځ�f$9��`�Jz˿�.3j��b��`z�	��^����Ќ�K�=�l�U^�|-�1;� 8ф
?r����������Z��.�����.�j)]�K!�x@�Nbx)0 �z�	̴\�v��C��H�i�'�\���Q�[믙:��:l�~�u�N:��g7܅���Μ�{N�9��QL��- WݢgR@�V�g����+@6~���2>�T��`��	R4�{#�J	� �~��B�8��_W�:H��j�{Nf��uH�x�� ��� ��n�CJ�'����$���1�i��#���_���x��d'�D-@z �7�Z���Έ��e8�O)�ӳ@8�&��{.�*�n�B�zGe�����z!����p3���s�msD��͆�p��=�i��Λ���%�5�\�	&ߠ��E-�(E��x��E[��>��u�Qo efB�������i+דek6��s�?'�ٽV Uh���4;����S�ư4���ya����md���¿4iL�`Kl|q��\1pCz�όN���D�~C���5SNxv�b�|{p�]<���vQ)N�z�8�Z�<Q�(JI��P�?�x�5dM/�Sj39�<�±d�����2�$^X~Z�,�����l����ꠤD��
k]/�*~���W��M�7��D��SS(���-�늪5ZQ�ʟ� a�1	��8��6�=�=�f��Ҷ� U{�V-�L��7��a֔&t,������ƒ]B��g�]w�P��i��{���z}��#
x�6���u�S;U?�p��
���m���R�鞌l�� ��jR�Dꇊa��QiR���Е��[�WR;j��"2JD�/)03r4|�T��#M+�>��
,�䵨l=NE�&�����i+�l Q�]�,���(�>[C=l�����³��)�H��/h�RI���꫆>2��6�zL6���k�p!y�%�nl"��8(J1�1#���v�wa?4| �X�&	�qŻ�Q5��i2�����#�-?�6�2+�g#�6�-E�P���I�e�ӴYv�d�ES.�*�H��g�TFeܷ�*TR��`��B����V&�#�&U����$��/c�$zC:����G�M�5|Ѿ�N����۫���2ۑ�:�.�$�:&�K�޹�����l^�����t���T)�\Jo~�wz�n	[݄� mA�
)���� ��%�������h�#�'ߗt̄Dȝ6�a�Y�/c��������;�+SJ�
��6��C/V;�%b��1�I3�+�;6�[��'5�%4��6>���(����+�i�*4�6�5cf⃼�jzq	�+䃶Q{���@�wH4�x�m^�׍F���.�,\�Ũ����P��
��D|0�O��*���ܝ�{{:J�?�ZA��5�g��Q����ѫ�J�C���Z�8�.�W<�5�4�;m_�P�U�����ds�gA��Y�s~�h"�G��L&o1��<:ڑ|Q?-�Kd�iR-��u�gڳ��㪔K�;��t$�����>!3��Ӏ�n�N��90\����������4���v�uٵ���w���4�T��Alec�����T8��8�j�� �w?7�{�HeF�!ɰ�����
��|�oD��N���r�}R���wI)�}�"3wyc��aF���9Y��V&=�<�
�͆����n-�=F����B�ݸ̬	쯘Y���Ʋ�R�wv��>T�n;c#��=.�ΗNh�m�cˠ��>:�j<�1���u|e%�Cu_�/�!5�?w?���
���T�ߍ٘%!�w�sD���M�^3%6-S�ݿ
(}�4��#�/���BL^��m)LOB'�ǧ��zh	�PH���
�����L޼1YG#��׃'u�q�-��
��if���lT�o���S��������8KVV0ב�!�)e�r��h}R���|�C�T�a���ak�s#����ޝn�y/*l���o�`6@�.�Fl�DRWh=����w���"n	�)\�^��@X���d8��Ғ:c��j.�J��|#�ׅ��AڞM����0q������=Iͺ3���M�������f�U�ZW��V/�ɏF]�$��gpE�1�a3�|�UF=/r���&���}�I�["/׮ż��+�&W�r�4����0��{�n�����pC�{�r�Ǐ���B���G�L;�{3�<c-;e�w�QeJjH���"���t�H��/��i��v��ݷJ"�;ԻgZg�ü��k�7�1���$�p�l�`����FY.7p�~�gZ^h*6;�e���Y�r�[jI��r/Y��#��B�R@v�	�	���+뻿h��>�h=>e�s����%z�s�N�f݃G]�LN0)����w�g�6�a�x�Z�A���Q�k�fé\S}3�pf����xk�b��`�~�K����CS0H��}mQ`��0}g���K?-�8��w���2@	`n�(��z:��$X�k�`�)]� D�� ��	�4��#U�:��c>Qe��7�ܢ�m@b���?kx�&�x����ɥ�ω����q���V���t���?��~~gj������i�%��>�Eᳯ�v�����$:��<U��-��eQ����S�rq�9��痛sIAֻ^�V%b=��Jk|5혞V!�w��o�gUgر��Pt����=��ڹqI�w�@��$_y�|᠟�i~5S�ƥ)��,��_V?����9Z-�H�������g��X�[G
����f'M�4�A�,eq1sN��nt[�h�3���m���(+a�F��9�I�:�*.4�/�����+�P�BIx�u8�$�Y��z��$����aU�0�=�h����{�"E^k������/]�c�X5�c)�f�|qf���K����>2ݏ*��;�;�I�E�,5��n�D�D�Ø���b�X�C4�q��!�1����.��5)����Mт�z�~��Ў��ʦ/��L��Λ�>5B:�h%�Z���^N�կ!�B�N{�)"�V��+~��-P`�N��?�\X��<��L�W+w����ڊ��j ��=C��3�;�N�+C�,ȅ�G�H��m��؍C�{�Uo�"�|.\�*���R���z��)�s�ttR��	�k�)Z�	�o[-,��\A��@���1�s�}��_W���If���Þj2�H3w�U|�8LIѻrr}�̪��B\��D�ڟ7o�N`-W����eA�H��:�t�6�J�v���	)
� OM�kY�N��νc�)�K�����.�H�ǟ�V|kg�b��U�%��؋�Q�I>��^-�|hQ#�M̶$1��?�1"ۃ�aSW�q$Is}��]���K�o��e����Lb�"L�~�٨h�nV�	H��v|C��ha��;4L��>��i�Ad�m�Z��G��Z����o�=�Ȭ�8$�Ѕ/�
�,�?��T�_��E�#�y�.�TN��R|x7<̐c>�j2Y�k]�4j��8�\��=d��䓟:8�K��7w�R
�ZB����/��`�x��^ك5��q����F���q@E�-+O7/ ���h�N��`�6���5��g�

�j�*�F�MLH���Y�a�����:�l���R���{Ԗ�L=;PZ�cݭ�9��$�:a�F�-���t�0�j.ƙp���[CR򱋞`����=��Te���[���V�,��	�����*z-0/�K����?6��.��;z�ON[0���4����J1�[aว[���R����1m]���H�������W���V�'��b�������أA����fC���ws��x]�b��hK���qZL��h��^�������'�fۼp�=��=� fh4�0q�uLCѾc8�G=�w���-�*i(���V���xV1ܟn(#I����L�| ����2C�)��b+��H�+l;DǗc�=
@f��Y}�a�t�~<�l�.�vo�`���5��9ڷ����~J�rj-��o-�v*�32��ԉu��c�4Gj�y\̔{XV���9yUMoo�^f��{�o/�hE���cH$��5��j�_ b��XSL7�pe�g�
̷
��c��'���m�e��	�ۮ/���؟��\1�T���TJ�<�Z��Sg	gy	���(0�Ԟˎϸ��f�� ��2����T��äꔺhׁ���,���g7����"���J��:�0 f3z��ߩ\���{fL�p09��rH��=��ʩA�.u���Y��p�݄Ub'�B�N�R�2��d:������hh�-s(-n:��f��p�#����[�q�Cb�$�%T�^�gQ��XeY蟳���U	�d��څD�������~��I9�ģ3�L�(-������o�5� �� 8/��!.qq�C�\agK�Z�Le4����{7j�w*]���[4-I��F<��幡\|�������c�j��/%���Ơ�S���7�����8�|f��d���"�X_'!�R��-�ý�K�h�Wݕv���`��s���ҥ��#Zm�$��_�ǩ����
�!p3�B����ς�#y�7��:w�F=�p�6:��4S9X9	�~�P���[%���dq�G�����^��w��>b[�"M�_
�{�K#��l=D����j�.�ԙ	?d�mHf�MY)a�0�kw����_��~�(�5h��M��7�j�n�Hz�nf`�:+wX�����O�)���HGH)�%����1ǒpS����]���J�)R!��ɯhG�$���G@uQ�wޞi6=zN����<��/n�")ЃpލEFzZp��n�A�7 �Ln>�����q����}����
 $P�(v[�@��it<t��cĕE��~�T>����-�䖍T`�c���:᝜��Ki*�^�@���~_^��ʍ0�S�/�Ib���2�aד1�~�F����ˤ�r#�"#�_@�/�aS V�����A_X9��}u<~[�����`���}�	�����!�0�|��B趦,\��9	P^�r܄�k�ϖ�c�fʀ��*!��7�x�O]n,�F�Mj����Ă�/1壋])̶��4��v�2���oDH���]>��{J�ّcǪ���m_8(������v[B��Q��*�l7j���ơb��v?�?���)����GRS���>ъ���CouLLk4}DH{�ZV����U�օ���I�"�-���+�E6-��ߚ���)�l=�'^���W,-�B��ic���e��>�`&u���A`B:�s%^�~y,�?d�m&��(����;�'�������@]��U�}f����z����:��Ɋp���ֵ�K�W9�����j��\uś�����m�k���S�H�6�o��[�6i��"�Y���q~�V(4���Α�]����4@[WL�R���&����`�A�^׀��pCKàB)p�T��ѥ�N�U����6g�p#��MӚ���ɫ��=��j�J�~��S����yP.]�2uI�'�h�N��Y��i���OA�Πk�����I^S*]��èA�?�-/���c�6^����>
AHŧo���>����Խ�N�Xwce��ޑ�@%pl7ڢ?6��'���'����������u+ԄJ��U�eŨ��|b>��m-o`���������93/��Y�/v�āH=׼��"]@H���z�L��iu�ԢZ�JD�~�n=�H+?ٹ���A1�T�:�rޚu�CQ�K����T��Sl��ߺJ��4F�OfƢ��C	����I��q�aZk�Y�`���@����_�R��o`�o�eN{c嶞F1;З��������ow3������c�/�2�ζ�W��*��*l��_�+Uywl�Z%�_h%�3ȇ���_s1A��mڃ��e*��k����K�Wю�1�xY#em��43Rw���M&6��Ցŷ_'o�)w�����a'����;I`�P2�&H"^Ҫ�o��#�}Ut��V�a_y��=��imGm�[h��)J|M9�b�AtH�Q@�e�	����
���+�a���	��>�@c��wd��VR�ӣ"����W|�YWC��
�^���'�S�(�g,�^#��|�� &_��JJP|���*EH���	�2Om$$F*Ab�H�����MA�q��$���U�;�Qr������Mzo����ޏ�QR�b#.�����6��T�B�|{�?W(���e
�=��-w&ߎ�7X��ng��QA���:\��эW��H�I�&Re��9�zS���u�����j.ځ+0�	�a\�/�<�7�ˌ_���P1��y�H�4�Ҙ��� H�1�f~j`/7����A *�@Ҳ��|�O��zMW�[u,Z_��������7�;U��_KH�#���޻	�o�;�R���ř�o������"J�_\f����-W���&^�*%�Ga�[����8�H47�f,%	���i�@z�~��r*<����۟X��.�<rlI����\͎�_x���_1i��T�Ehɮ�KWI�CkO�H�=��4�$���:E7>���A�'� �RD��<���Cʱs��^�e��Ĕ Z�e��?zE��U��qs�?�^Xg䮪? �\���7�ty��9HU�٤�6:JeGV�;��Y�N3R!R����pL��.մ_2)L��T�_D�Ra��~�����P=���|X/׼��}-����PZ�w]��[�u8q ����	W#$�˘I�y��?,in�/O�ݔ9�ccC�5aaj+l̼�����H=��0~��$e����F�0�t$j��`T�*�ug~\����T@a�&^zJ�\�W���;�M��@����g�4�;	Y0�R��C8��X^+�Ugsv��}��D�zC���!��NOEW�.�Q�_+aה/"ۡ��ި(1BʼQ�*�"��\&����=���W�\�A�bP���*�?�iI�����a#U�YB��շ�7Rϟס�#jr�f/8��bfؑ��hٚ�P)g[a���!�P���Z%�������I'Ph�ln���}P7s��{7V�y�aT���#5�2��oB�Qu��v�����F[���v��*����0������ח�$Ef&!`�i�rI�%h�廍�˗�O�dH�E��R#A9_U^���g+JHL���P�e�̖�>�ȁQ�f�}��L,f0Z;1-�./9�D]�Kɳ������Հ�JȐ��v�̙�U�[�,e����$��^��F�g�H�d%�/8q%dRr_���Pxd�/U��Ӝ��L+�c��͝���~y�0��$��[�Q��˯��E�Ϡk�8>i�����ٴH�{�Ջ�[-�jۭ):���(��:0,H��@��&�訫�W��[x�V�.�����(��U6���� �
D�{�o*%Pҩ7��F]Z%|'$��_&��y֐�l$��xD8�蟓����������6~��Y���>����F��G
X?j�ܲCU��z|Z^G|)�2 �t��Z6��K�&���آ)���2.`�>��Ü��S�E�� u0�I�l}i^iѐ����֎d9��r��E��/������ʛ`��l%��-��p��}�ʵ	��Wr��w�1{��A��7�Fo�U�����I�U�[����8XH��f[a��A����Ҥ�n�s#Yً0㲻�t�������&`A�bd���j���y['ӝM|�E�]^RI��[��m^-�Ҽ>Yp��.��4ABX��.��&���M>v�p����$��0彭jZ&RWԉ�5��b�q�ɖ�����
�HXN%Tƌ�0�K��/������� q4(>s�\�o��;6bA��+"À~Ԏ���u���w�I��^����4�MFY��b��Y�p�$T�ZB�uoO:j
&�@u�.V�`T�!�����>?���F(��t�g��s�}����c��[�<8�[�?WIվv�B���PE��� ����O�-w��{D�d.	՘����um�[}ў"2d=���=3��1�[05X���.���V�z1�+>��^{�/���M(p|�H Vc���SRSsY|�ڐ�5䗦f��R�K)�a���S5��M��rS�0����NU@;�zf�"�d=<�˕�t�7��/p���]4[��?O7�g�/�+�NP#M��m�E��s����t�݋�1U�h5[��[�0U��=��J76,+.۪����F E�t��ON~8�Y�n�Cx��k6��F��R�Q����B��`�J}�o�A���"��ҿ����x�J�.����8m�S7�V9�	(5�6���WSEGo�̮'��~������Kq`����uCe�Ui�#ٶ?��t>-[�Po�^e��,[h�	�ժ7��JPq���[=V���|Qje�v�J.>�!,�6��A�|����򪳗�BJ�Mٹp"H�	��t
$������HFpvo$�O彋��C�(&�ʢ�J �a\��n����w��؎tw��.ZR�q������f'�?��zz�;�E��h%�C���S��0�l��b�O�[6R���0��N`�Mt��;�U���k=+�2�ᐛf#�v,�U0v�!��8|C������ч��DL��j���ϗs��^Lp"?�x!x4�LSV4�6�l�4i���UW>v��rO�{@9��:L���&a�����\mBHn�����:���h�v��5e�fG:n_|SV�Ԃ��*����HeF��3����䞺9is^��q����p�h�e���XG��o�}cO��1\�&��|?7{�p�,��u�R���m�� X�(m��ɥ�G�����j��_����["��}I�����'�E�I�p�6���Ի�>(	k�'?�b��`}#QG�#��w�� ���)D��;�c�_���wꂚ���`�#��JcYuDyp�~��B@�ڑ�&6�B��������pg�^���#6J��R�8d��My��v?�[ӄ_�T�����![^��J"χ ������{�XMN0�Y�������`L���ʲ�:������
�����A�;���Jqkq)Z����C��)V\���n��ݭ0� �о���g�b����>{����$1��߇,(�Z������ w��t4<�g��]�fnt�^�}ͺ���֚���l�����A��ݼ}���$
��|�=��I�ȵ��_xQ���WUם��)؉:��6ʳ�¥��t�(3h��V�֧����{Rz��9�nj%�� �ٍ/y2[ �l�v$�]t����U�9i
~Hz�S�MǏ;v���}5��j�5���Ɠ��w[a��� A�b��v���ʹ���5}��i����3sg��Q�i�Ea3�<f��G
x���KR�uY��n���uo��3��F�d'q�)d�r���}��v�SQ����Q�ߪ� ڿ��Oa �/ؤ3`�~�P�1�4��ʮ�����L
)��=x��.�-��tj���_���k~W�T�y��i��u�ܥe��i���]�����4��=Q ��M(޾��q^�j�(�G��hc��M�yq���Ԣ���|��]����D"���F!��5�ss��*���[]���+N�jhZ�{�̰��|L�؁��/t���8�F�k���n�z��x�g\��q�n��d�h�nP��� �׶�vy̳��[~r|w��̟m�2H��ϏI���I9�V�
�o"ih�D��:s�7�9�[��@��a7��R�=6��ʸne�?�I�+���Ѹ�v�Jsw��Ie�I��axe�uN���O�Q.ڱ.�����;H+n;��ޠw�Km>#*��Ibl�n��tHm�]ޢ_����ImE-�,&�T�A���ӛ���ׯZm%@)��۵�T2¤"/�PzCA��T�J����v?�>��#D���*z1?o�Y.���Ш1m�a	��H��DðE��}��FX�ο�|80=lck3	�L���Z��;kl0њ��O�%����{��(�p9�[0\���R�	���9(GK��y9�}qE?- ��3P�.<i�zb�e���d��@(2� ���Tt�W� �	�����5mm�Fr��a�<.��p7�������g����qg�˼��Z.���,��m���nd8�Z
l4�_��5���_ _� ����֙8h򫯖��\)�6�/\�>�b:����..W���ҖY��c/��n���mާ2�Bt5k�g�|Zg4/x?�7KC�כYp+��H�� �vv¾$N��������7���T)
���`0�����k%���vK�%���>r�ѳ�FG�l;�[X���~���3��t��1���u�6��B ��G�o;R� ������'�����VU{��5�N����.�q�%Kp�Ř�E]�~.��g@�%�}0y�s��%u��Y��kͮҥCn�;��ǭ��P$9R�������d�� D_*vV.��JHOO�ۡ	�������ؼp�q����?���bP=��R�D�$Q�>M �j	���[豼�S)�7�S@c��! s�zc�㚪xƘ�Øg����a�ɢb������9MϮ����l!��]�p�쀋����O�2��ŧ�B�a�w;��F�alޤI��zFg���S�4�Qe��{�����-!�A�x��)��u_��G>���%��mlNDoe)6��:�'z�4�Յ���XR�=94��,��<>���lI\2�3xv�r�Z�h[k�M��i����{��WL�7qڼ�z\�"şz����z!�� U�7��I�ͼ��e�5m��b6r&���}ln�=u|����,D����4��"D��|m���֗j����G�M�:"���$vyvze�B�U1ֵ�O�wh�X��z���*��vN�^"��1���������U��٨f��,�iL�a����A�OL@��ž\H�e9i�VP��h_�4܍�$*�h@G��"��Ӯ�W}����@�̉|����>3Z|S^d�&��K���:� �쯁��=Z�4���� �K��@"eo�����E �nA���B����F@O|�K4c{�C�|b��O��3� �t�h9�׼PUt�|���r5%j��T��00[Oƚ@����j���U���4�T�&E��!3T25Q�X���ܻ��<�]./�)��oQ��_%����C>TytLaW�y���8��W��9����X���F��A��k���[�X�8�X��'�Ƹ�&���H��ú��a�o�h;p�5��{3�eb<pe�0I���S	t��6NJ��Z�-³��z��/z��g�9�ďEh��:�@���O�;GڕL묟3(� ��f��/Ye���z��>���f��k�/�^}�î�̏��~�����Du��b����P�В�6<>��ٵ��}���r�ܥ�_	I�y���M%�6������Ke7����,�I���r^��1O
B��t>�Z$�QW"C����W)�ƅt`U.���/ۭ���lG}[|fؠ�/�G���vd�����L�6��7�y���Z�C��]���>�P\�3)�L?�H�Q[�<n��}Hb-f�?��Am�DZ\��66	� 7wW!�;M�����r��/˓d��^��#q���F&1�*��jښ�W�K��dh����MT�j��Fp)*&��Wp����O�N?X��E�lKN���#RmDF(e���O�gAi�����:6���r���:z�O<�Z1LY�᫕�u:�ʛ�F]tc:�B"��?����V�L�:�݌������H��z"�������"��s�J�Ĳ�-A��X�N�Қ���5mHy"�=i�0k��T����n���숀�������[k��#�n��43C�|�/���e	�֬~����3l�VphY՞`c���"x��P,�^�g��l�������� VP��Owa�k�p�Wh	_�=kz/s{�,D��<���۾r��)�����1�]=�{�춚�|�Tm9!��=��搇�<�f%���U\%}N�Syn������cRK?q�c8>�T�uG��.�β�Qo$�6w�9S�ДJa�Rӂօ6:������۫I��Un�R�������m����P��V�G��0��g7~������o��h@lG��V���&�N�a���ԥ>Os��&�%z�hV;KBɭ;K��gߋ�=�4o9Uэ����ݶ�G����m��
�g�
쟍�z����#�W�m��� �}tR�������~t
�KI���� �8y��x��d/��]GB�������j�c��NW��"F�O$G��R���|	"��y�~�g�x_w���ڌ5�9M�R�:��ێUj1��嘕����������(�4N|�;Wpi~���v�ؕ����fw����r!�	P,S/
}c�^��m3: �#jbL��CH[k\�����Fvr~J�r�<�8qp��4��ĕr���F���\�:��b�&��m���qm*��-�-��k|7)/��5|C!��Fy��� �~�A�vk���{>�z�ѐ�;�Q�Q�F��T@���yI�J���*�VU���1�@\��(hi&O�W^b+4���|��E�Q��s��eQs�d�n���uk.p랁�! ��ft:P�@�m<Ɖm�d+W���|k��(4�4<g�K?]��-���oSq��[H!�R�SXC��F[W� �w��H��e=�!���KJ.%S�;qu�7�����E(���WB ��w�u}f5���
�3�t������Ck�sxȐB��Tf�#q�_�xj/-�K��m @t���@	DwJh��ű���f\(�ۙw)cG�sE����X�I���hF�ڿp��Gɠ?G����r��"Md�P�fσ�I��t�Rem!����2˼<#�:��lX�Oo�_���@G?%�[TC(�t��-����O�]�qB�J���_OC{n�EUr��zDP	o����x�	�<7���ÿrm��|�����:�+�D��$�������CH!�����(��W�����3�g��_;]ԍo�kN^��W��/�>��]�Ě�w{r-d�ކ�I�`(�� >?M3l�R��V�)t |S�poq�&5���o|^��Hf�zt������Ƹ!��:\��.�mez]�O�ՉǮ`�^.,�f�ʗ����3V"�G	�{���n��S��	�ᇤ>}��_�s�ݐ��B�1"�v��J_�x
뉦w0pv���o]y�M�.	��"+�п��}��O��?w���^�����`_S���Z+�7~4(A���$9��O������sݸiX�甈CM�i&dCĝo��g�^yu �cWpq(��M�+��׿,����w]�r�/���7|��^V��"g*�:�|[ˢ���Œ��;!�ˬ2��x4J�G3=�2J\�\��N(��o�?G�ӈ.к������hf�n���Ay���y�+s���aU�l��解6i֛Xe\jK`Er�Eg�Pž�-۶��R.���o[���r�����w}�Y��9�WG�c� �0rI������8n�S�Қ���|��s���qk�`!1�B���:\ܲh�2K�_ֻ�(�&&[d�x񶈔�L�K��&a>����+O���X�������K�����u��`ɩ� #�FN>�'�Q�ͨ+ ᄘn�6��m�W�e]�.�����'��٠<v�_O���UFޘ5G��bo��D��V��Fg���<Ta�lv�C��\#�n�����V��s���V��짨A�.(�����o�.G�*����j���z�A��9��8�Y�0쐗���-�]��<�Y���tC~��E�8ޜ~e�������'�J�3����y5�P�����rR^N���ٵ	5�x�]�U���=����_����� D���o�#\��,�(�r[6�=c*;�(*��R<�o�F��W�m�}r)��i����E�ޙ1��/�����:���T��n���y���l�,�pQR&c:<���@�8CfG4k���Э��j_hf}�v"Z�T�M��~AQhig��yBb��Tq�S�ί�/�m4�"h�=�v��#�d�+�[D̶�W�N�oe=��>]�T��Xc;�;��0�n�_;���V��G��n-Gyڎ�)O����V?�R��2{�:]���;�S�D������B���c��T慯:7L�bq7�}�̟m�n�?U�þ[ʓ�
;�D_�p{��y��?��`Z��,��a+�ם���zؑK��XM���[=���aͰ�+��j����}Ο���V"\)'q�dw��!��5-���5���W\}���QD��ƟqqQ��OϢ�<@P�B�!���n��¼x�/�m�&���F�2MW'Ts_X]�d!�j��a�V�W*B�C�G�Y��lx�0�J�V��ܥf�0bw�:�8��N��C`ג~����i��b�H&J�������� V�ǟ��v�k�[C�{��a0]�P[�� �|r����B��u
���xiW[޼^6c�33�X�QfVKg��l�u#�Q�[��԰i�S��0>z"�{E�l�l�8ȥp�x��,<4�,�:e;&ޕ۟6
,�8�`�\Y\�p�涟��7xK��
ycq1W.�hJ�o�M�0p$�F��	9�qI*�|� �<��A��]}{W�޸w��V�uwg����o���t����]ZZw�|&���6���	��>j�+����rp?�۟�g@���g�@{!Z6�@=��[ע����q1q�z�7�gg4��Ϛ
��3����T���6�����o���ɑ���n<2҂��i����䘖�$L��q4��ژD�l�k��X���Է�]�ϩъ��.�-N�N+l|9{M]ZH,ҍ{��E��Q�۸�
��j����N���Y���,:��$Cl^����cq�<tX��僽�J��;*�>㵩��|�Xan�J��:o0���D��}���Ě�t!�cSw�������-<���2JǧQL"��-�X�P��R/�qWQmo�Ph������N�7/
��tI�0�#����	hy�D^�����w"�ӝ�:���[�{X�@P �����X8�9��܎ٞD� �F� QGs�x�Q��*����|���(5���k#mfש�"���ic
\�/\&7_O-S[�h�Tg�׵ח�gRn��_8`��X^�u�a��݉���gszNk�1�J����ƇY~�Y�:e���ia���b�� Pzxih���;��͢{�4���N���������M��Ts����8�e�z�����[���18dfӋ<%��N]�sLPG��X��6,���4��X��!:{ꈋ�(#Z����Cg��}壣<ʿ�	t��O}����[�?#`)�z�I���۶X������N�llB!{ȩB3�x�L��>> �4��r�q6�ARE��V�	�b=\<Y�*_�Y�\=v8�~(�����jF,�0{{&�ظ�bd��|h��a��W|�O�anT���hLwXϢa��*��$9g�[^���LE+mP J�[k/Nݴ{���~R���ج�+2��@o=�	"��y2��).}�0������.ۨl��<�mM��KA�����^?�0\}!^�\B��#_��D�B�7����<�E@���pG��8�:�Y�~^���g�񟪇'ϵ��.` �)��ND�f��V�¹�e.!�� �sE�"�W0V��zf;�����C�����X]��g�"�ؐ
]�=<�j�6n�a�[���K�ڳچX����Ճ6��sb^�Ү؆T��C(�ש#Z�	��e����({D���Ž�hg	\n�ٺ,a$�L���[�����+���:�:g�m��\���|ս���Z ��9L���e�`�T����Q��d�����.����w�&�R0�Ȑ�Gycu~�t�w	 >��Z���z�nᏒ���?����Ԙ��Q�d~�J�af�'�OY1mկc��2��V�Ow��eJ��M�Z��E�8������c!pum�R$㓛�jWok%%�����6���_�r\�����Lp�|�u��SÚ�=F�6r�y0��,0�����a���qS��eR�݊w��u�&h�gf�g�V����"�a�OA��:ؽ��w�&�͕�#�[&Y �&7�����Y�-K�v��k>�_�:A���k�*�c���vS�i�������wf��w�9τ���ۏ9w#ok
R�򽴞��e�&�MY�G��[��[���Ew��O�U�&�h�e=����
j����R�~�n_M	��VR���]I��,a�f�N���_���jv2浗��g6�s�4�km��g�?��"
4c>�����1��5ݿ�R����h/��������{�����6�rF�|�/���[�;���l;�^�����˝�i�5a��D/���1�;ל�c�}���ڀ;Դ�(q4GeU�y?t�x�-So��/���؛Q?���z�-����^��s�*�1�Ɇ_�Un��(���S���!�;	��Ţ��d(r(���[�ӷ�p������)iXg���=)���R��v�G}��i,ܼvm���gv��~�G�0��(���n�`n!,�dԈ���eu�g�= ��CN���}&>#��1�'�����߸f9W�ђ�U�%�Vgfkod��q ��M�7�'���sRB��fX�����F����6��m��qw�Pdlb.~a�eq���Ʊ�#X �a�o8~h[%��J})���"vxI_�
�1 0�dK�'T�j�k�Jy�mƬ˫��I��!hٜn�v�6�7�z��>�xR�G�k��h��26�q&~���m�w
����Ĳ�`�` �9�m�� ��Irwx���J�t�����ޛ#c�i-lh\��`��sF�j}� �pY��&�������0�^��uσ��{�2T�Bl$V�q���m�Y�r���c�2}��P?��mlI5�|�樳�0���>!߽�}�۠f�d��hl[W�˷�"Qi<�N����6~������0/������JD�J�a���� �� ��!ٕ��(������ד�Wi�ܨ�˵6����P��J�V�j���m��w��X*�&Xu@[v���ӆ���{�2g8�e���s�y[�5�d�3��������cX�Y��e%r�]�j�ϔ���śS���E{
�m2rym-,��J<	�!�C���Y� g�x��8�Q_'"$���������O�^6��sQf��}�@PP�*�!�����n�Xs��ե8b3֕�e��܍�%P��C�&]�����܀TS���?y9P	������p&N:��eWq�1���8��Om�v�&J4�⇅%��@B^���Q��+�ϩ���kj�?O�����-/��ٷ?ɐ��=P�l:��g���x��P�?e�ܦ����B�����O��������OA��@�]]���_c���X��N��J'V�UV8�05��%F�6�׃�.{�|^o��-\��h�xP�n�+��AG!����4��yY~�}��i㖗��4�<�箟�"���8�(�eh�`��V�0�㌥O�c�h(	:�%����l`4D;V��G/6 BJba�+=��ȍ��ˀM:s��ۊ����x�@������ꁢ�$.��l��A6R*�C�x�ɥ����C:8�I&��9t�	��y\з��������tk=%2���cR.�0�����q�$hј����wO�.��xpn3t���p�����lz�G"�߾�ݱ��?�1��+�k�緢	���kr��}�%d�w��'�H����d�u)�:u��*+����j�өu�!��DU�T���Rrr�U���q;V��i��4��e�	��"��g\�Ȩ:S�a�X�Bc֛<����kx[kKM�`x�Rv˓�6���&c�_�-"&���p�w�v���<��*k)�IP���S��''{%��)�yh�DΓ�ry�p�GSIU+f��_�Xn-Jʘ�b������%R�!]9���WJ��X���(��I+�`/��3�����"��\C@��9�9�*.}��cy���Z�|A����xF*(۲b��0R������ǞF��p��;A���}�����A*��Y�-"HU8
���`ދ����9u|� �S=A���!�
��=X�)W@�*,��sW�Ne���1
�>c������"��#�x�P��:ir���y{n�D=i����Y���G�+�{}{֕�d�H�V�9>�׼��� \�8��͟��� ?���~ѡ���x�k��4����7���ynD�O &��é@�#	f���ܩu\����!ys۟|g�e�Կ����v�+����g�f������x��X�t{ls�$R���$0;b,���l
���Q�u�@L�{60�[.5a�7�L<=�E�T���s�>��;�C��0��;�k��:�G"��T����gd>���Ą"u%��LSL�)��#�����~K^b^�3�
�*�,^�q����hE��������Ǿ� ΂%�%�Z�Ϝ��ąyu���0'YO���s����"�5�G���|#���.(���k�`bJ�c��HTEk�EN�JW�Z��U'�����+�v,�m�NWx�q���̴�V�F+���H"�h�{^�R6t�H�rW��K��1zҖ�_�׿&Sv�Dt��J�����T ]�c�UN��.���G=�O������&���Xb��l�Q�a�q2m���zrB~��Ұ��S�B�u��fݯ��L��4��K��y]���iEl���~z;Mo����;�E��$�x�[�ײ]�W���� �3,{�| 2x:+]���k��'���)���b�P\��w�vG��*BVzJ �Y�ԅ\7�:X�>�z}�_�[���AF�Fvs�\@&�7Q�H���t���m�%�PH��v���!D�(�@��O�h>o�>�zQ����	HX]M%���q��Ը��S>��5�Y:�
��	ӕ�@�
W~%2���m�ܝ=�'��F8bE3@t3��n2��)��@»f*9��l�.2���wH�I�$���ý�0�����5���l��л�k��֐.J^?l�ozoVr0��C��	�%7$�H����s�K^��t��5I��
6�G���7���nI�������;?�7j$�-p!�[q�˱X:9���d�R�ٱجZ�.���0Y�.�f���ki�T�* ՚;�nj9q�MXQ���;R#�2�:�
�*)$�Vx��
��]�BR,s@�Z��a/;�Co�����_;����
�o0>%��'���Lm� �c�xV���W>����%�c/
�������^��g�՟�J[�������{��sX�x����b��i�T���䢇JaE�E��h|��N�h}�xtf��PR,��P�S�~�c��U�/�p1[���\�S^6T��2��~��B��Rˬ�Y�훈���U!'�'!��n`w�f�G�s���tH�a�{�Y���x���÷�ꞈb=XMS9�o�(ėM)�ԓcE�ּk�i`HA��^��#"}�Q [8���>���w��Oh�R��f<Y��e��eC7�8�fb�37��vBh@l��HܣoQ)��*�r���}��U�X?Ne/�(u��,=�h��̖44���=�.:>�}�gu��Ik(��[n����k����^�՞�"ņ)C��`�B��AA`Xz"㧒����+{���������p<�
%��u\{k(m.M��Ȗ�NE��>�r��\%�:o��Mp0�hJ����r
Uf�|�� �sOF��ci�C"7��
?�_�QR��,-ʙ3�|��"��J���,��ϐ*��N2o� ox�">��-{Լ+�0�:����l%;������j�����A�+�13:���*�;��� f��� x	���*P;uj����b`j�O��u-�� ����������YC08|qߜ����a�z�fS4L�Rh�&B�����U~'2r��+� ޿��ny%#~ܟ׌R6�S���=��d�ѹ�*��s�y]����r�]4�`�$Q���Kp���q��G��VxEf�k�pq|�N��]���<q#�j�/*j�e� �1��q��[�p�5VF�Oaf�����]�*2�A���iƴ�x�&Ɣ��C�������r0��a=����~���/��͢G~ /|���{��f���"  C1��O0}����4R�z=��g<M+\kA?�][#S���r�e`�h(��"N@����E�iq�;���vk	�O��'rWZ?3����f��?��!K��}��a���?��{w�UیF�������#�WO�kV��4���܇>�p�	���q��]2��1�I�ZQ���D��jRJz�]z��������e��E�{�9�����I�R�e�b]�Fh�'4ig�5�������(�8E~�me�o		�"!^Is�y��0�H0�\q�2�}w�r5��о�-?X�\�b�M����f��j�����4�kb��-=wE���~��$ͪF��܃\��h�l/J�ؿ�b�ߐ�J'�@�~T�?_n�F��
� !�SP����IT��1B�,�9�[�%�?7;t������nL[Y�D�	���/���!�&�i%��9)0&�;:�ix�lqc�o?�B��(��f^�H W��/���f�E���~�/�,��;h���:ևE��o#���o8E��3��H,b_�맯��;羦�=���[��ܞ�')�6���g�s���ڻ��C9�x��nz4�2v�ڐ$�fqe�e��F���X�В7.��.2_�(���KL���M&!�OQ��)N7d������<[�?�+"�d��z]�>��LC�U��BĈ$��/�<	��2og2A�`)�H��������hw�0��y�G��Hʩ|I�ul� �ƿ�DC@Fl�c��!Yh1������3磡2�ǚ?��G��PT���>fW���c)���~�z�b��A_�Oԅۢ�%)�� F�]�	������o��g��K��Ѐ+�A�
�E��k��Z�a�kL�P��D�!N΁:$���f k�<��bn�_�P;�p��!&<`)E��Q�
&�t
s2�2$����fJt8=s��r!.&��N/x�".s*;�˓�#���)�rp����۳$9-$\Je�L�9�XU
�b3� � +`��G�·7 �(W��҅�/�T��gu���̘���fJ+�_�,p!�/�|?�ݣ,���?���_W���ٵ�fet�D�5U+.��Duy�Ñԅ!���:�^&� M��F.ԃ�M�UB��a��X�-�������IL<�O��Oso���b�JVĢ \�/&?}�kt�Y��{��� $�].�6RnF���#��;h���s��m���F2?5[.S%ڂ�����i~��G��˕`�}`'����l�Y(-�M�0��9�9ȋ�4^%���!�x���C��H9��X3,l�KK�[kP2DT)�PcN��l��\^U{WF�5P1�DL���s�TA�� ��n�|����������7K�(�+G^�2_Z�����Z%����̆⃱x�~�ggbVd���җ��|��x/7��>r*j��|�d:P�K1\����rI����]'��0�{ٗ�~R�G�)5�B��炯P\�2��Q��`D!�"2�{"^��ؠ;Yh�@Un�3��&AE�ߗ÷�-�Mb�>�G�ي�hG�p�	ba���ꥡ�K��Y��pZ������΋k��p����� �x���&:
��`5���C$S�e�Wn;9#�$�$$�(��G�u*��j��a�}�$O��c"��=�A��I�=��q �X':8)�%�_i*���$6���lB�/�d^|k���|*bït��hx�J�:_A\U�PP�����z��4e�Ƞ��T�5��r6���Z���ml�`�Jd��&�>��ȍ�����]�l��S��ץ���9�����vb��o/WI��p�_�5��(�l�'{�?�I�5�l1��y�maK-d؜�r�Lۣ�E�����ʳ�(\��d������4,J�#�V�6��ԫ�B]�x�D|���_��^$���.���bb6�x�b�vc%���!�8�"�h�B�f�vi�}5�L�����;��{�g��v���X��cw2�k.�%{!�^ ��s�v��d.�_�~MQ�k�y���N�����;5����u�� ��
�'^�d\Z��U���G�?A�)
���C��@�V�ޙy撌�aE�="T��1�<�/�����e,{Q1�7_I��'+JM�z�MM<Q�u���Y[	�n��v�+��a�v�7��i��f-jEwe�X��{���N�:3N�B�{���R�����3���:23�?�kG�#���ҫ�j`[��e�Y��,/�����z-�P�e���1yk�;�'qw�3�����,@����������/��XgIp�[�3��|��	����_��0��P�;���;x�$GGXq.���(>�K��x� �~N(��R:x����IR;��ѮF�=��qQ�(O}f\-��w��O��s���ת�1Kۊ�l��[�z�ne�f������w�tt%CgH��2�ę��y=V;Y"���,$r�Q���f/^?���hL�7ni��o�(�75�,w�d���Y����/�Uv	L&�U�3���6�	/��F>����|O�+[;��z4�u>ɴ�5����W!̍�@
_���E���{��jt���g6L�u˓Z����\��Nt��_Q��nUe#�^�q��<9D�5�ד���%-[�\�9��Dk$�m��K�:)M_[%vj��Ĺ�K)������$}�S%VIE�BtM7����\P���,���k��1��N'���Ou}1$8�xT�����?�ӊ�ʷ�Y��v�f���'A�m�3��`0O�O�F7�J��6���~�'.����ɽ�I�4^�u;o��U��-�?m�����~�l���ʟLq��5��2���O�O���6�N�>G�C���Rd�Z��X۹��oC�j���ϳyL��b�d�]�y����c߷G�[��T�(ߔ�j��,uw n��~Y~zЎj�5��`H����{@.*�?~��F����s��������`0�Y��>t�E��+�4�Q�Q_�1w�e��9�VK�U8��\�ɫ����8ٞ��wl�G6S��\ת��]M��9���ߍ`wV��@b7cڹ��9������D^m��r4 D������m]!�r�P}��ŋ���rA��7�����7�f  @����?����X&1c����nC+��i���~Wz�p�I��Q�ٖ䈈Ė���ѯ�#7�����}u�����[+�����T��:N2ު
���SP� 	u����K��4������Dt.� �����F##�6��]�e_g<�@�-^��������+7�F��ނ�����&ks^=�H�*#YYj����5/n�^|�C�X�&/$��6T���M׈�]N�	���g	 ��x�c��M��a)�ԣf��� S$�m=�s�"���;��2��C[:_xi�[����@��R]��@1�牟|%Q�;�v����+�@�[S��0E�����NAwˑ�"J%���J��l,r�E}�2�N��J��p���y?�-ہ>{$��s��%>5Q�?���:`bOV֮nOi����������g��^�X������!�P8�BaE[/i��r�:џY[�E�	q�v\����t0���8�1D@��`�Gc����X;���*���X����=n\�\5zBEG^ ,y{������G.���*k��A����q��*�<B#�V�����El����N@��l���
X7�m��l~5=������?���6JoMwD�X�{�@��P �2#�n���]U|3���q��t����,��%�s�	��گn�=�1�	sI�xnG�x����t�jG���J��f��p������smi-��z(�X�����z�L@ݡ��M����ܕO��T�!\0Y��̉X����	)H��r>�����e��^��U5L�q��m�J��A����h�� F#)����'�p-&��:^�#����2�4O�	�;������T)C��G�S����845/U*ze���i"1=��ʺh1$e�\�t�_�_�&�+�/5
2��N���k!��Ǘq�8�ω;��loa���%�k�W$Ole�r���̢[%zJ���&�{����s������{����3�+�yxB1̺��"�:�4F����������'�Q������-﵍�N~���o����Z�8+����Lc�$�à��jH��z�_<<�#�4�����1��E�uҨ�1��%�����]��~��񫲘�e���[7HU2��ɫ���е�Q�ʫ��RԪ�]�o|����a���K���w�4�����>�JX�*�f �4�m�ԥc�	�U������B�1�]\[���>���s��2w��u�Cv�����ͺ����|5y��T�io��G{�Z�\�����N*'�w�3��j���8�Fۆ�8�	���a��P�f&�LW��=k��q_�N�.]i����S��[�Dv���%Kl���H[��b�:��z(p��F&�q�{蓄�bu�r�� �̌�w�fyZ���X���`����F����tbzD瑕��d%���r���<`���I�/Eު�m�& �]��qr�3M�� K�Vҙ� �DF!��$�o��Ё&~�P���D��[b�8~���C/��Lw��س��7�,`��kW���3����7�jW_(4\B�@$;Q� ��¿	���V-s��~Z��H�Z�4�aqX|�M�{��hb,׈�]�7�}�a~�	�8�C�QXl{���ڜ�0���� Ŵ:�[s�  ��J��S���?"_i�o��"�n"n�Z/�k�s���D4�w�<6�LҪ�w\�Pn�uOcA��2N�*�\����o�}W������\�s�l����f��o�Pp�ңh�'B�����c���LT��NE::�,H2V�U�-��'E�U/��][a+�"K�����Ρ��LL[+��և����$�tޜ-�'FzX��C��h��~�!�6��K���$�m�H�Ĥr蚇v5E]��X������
�o� �0nͫA�ïb��j�1/� �'�ٽ&H]��0,ղ[���DpF�����v�#mC4�kO9���p_go�po��%�?%�^�8F�M� ��?>������ˊO}Y�%o,�g��0��x��+xy�a#8�vzc)�s1sc��N���T9�ϯã�@�0Q;f[G���&��s�)��F鹝�Q^m+�u���^3����PIM\yJ���L,��ȅ�a�{;÷'���|f�ݦ����V�Z������j�3*��q|�o=��q���\Ƙ�J@!�����L��sGuwIإ����$�[>�ϐ�nϜ͙7>��C�"[�^��<:�SAv3��"����Ιh�mf-��˂��p��`�o���ⶆ]$G=<��}޲Z��y;ձ��?f޺+�������۠�!H���!hp���� 	������=��������˚��?��]]�kW����I�|v7U{ԥ�k[ZK'�8�B�;;�wh���Xg
iBi��)�ϗn��]P�!?��I���^�&(A�`�/+������7
��r($���0Om��ܩS� '���F>���?�q�Q�����#d��Ld�NU�N?��yx��4�����H�����^<_��#Zt�}詻����aG��]M���R�i���~L�KD�(CU�j/�ЕYi�����m^�e�����uI��#��yj�
e0��ţ��iFh����ӑW��������"̌(�����-l�z���U�x���I��O��@�F��*�&��O:�z�$\�C��֥X;D$���N
hU��Ө�0�*��	.bw�Y)�o��*Qz��n��� �~��E.o
i�;��2��6s��|����j�tłf> =�׽�ƞ�Ml�Kd/t�9�O�ȳ�ݯs�9}K�O�jL���K���4���ۯ'�J�[V��v�o`{�D�*�1g'�)�,hC^
B�ɯ�D"5?J��_��ד!��K(ij.l{�o
�����<�[�ө�gUB0��;��-��
����5+w'�S���,0/�z����T�]�EQ��c�N��4��?q�(ڊ��'�pDZy/;�Z����7.��,ſ�� PZ��oe���6�Nϔ��	�s6j��JK$S��0�&j;�e����/��/��\n	J����t>İӥ�542ĺ�,�[�M�i�f�s�oz��0����P�_ݛ�[�C`
F���a����!kY�����W6"��.K}U��ݳd��eQ�W"�g�����Or�Do;��񴠍����o'��ե���J���U�:�S��9���o:O�J�NM���h�ݙ��;P���v�ד��j���vW�~�\Ax�q
qk,�6R��#���+8�Y3̓	~+M'yY"�5D q(a���r�ږ�o�6l��qq))�����l�!����Lwy�Lq��Wȡ��fo�RQ3���K@���C�nq���C�PД���'�ʬ&�ڗ�FV��!�y�.\Ώ͸�(66�a�+3��gYp/���{�!,FC�d��\��10�R!+2�mp���I�|�&�xhk���Mu�`՜��{�X�٥ra#٤zL�ۇ
��r5���;c9d|�5A����b$�WU�"Nu)��Gm�]�iy��Vl�N���s�=-�į�]������K�_$
�z!� 3<��%k=w��W��IJ��+�F�t�[�5`�]�%�82\�	�9*i�I�K�}�|���^SI������T?_C�@��r3��vY��n�1勵�JW�Ib������!!Z�������:��;8`��h11:���LC
�������������<�
,��^�7�mjS�'��8A��;���^��no�Y�� UQ_��� ���������&w)|��6�y�m\�tl���B�Hi0w��\�� R!4T9j�������%�������Y|��贞[I%+o��}��	�t �
�I�x	�:'(k`�kЌ;�1��X(�`�k+�&�:<$�D�0ii����6��n[��+�eY�P{�':�����]|y���>[�hT�}O	����U��48�r
+{r:\A�éq�z�������.u3i򣄺+�iA7iʔr�C1�b�Xk��P��a����(."!��J��7��\/���xjF�����V���k�l��YK)>���5��`+NR'ǯ�D�P?��e��]5��9���s�x�9�Bƭ-�&�Рk�����eg��"!�O�??��[0�hz�I�S|��P�z�%�`��2A�Pm�r:�K��J�dyg�;sR@{������ ��������U�Ϫ��$K�������)EhƁ�N��w]�ud�WS��6b�_�"ƀ���;p��}b��4�ٻ��hf��sC�>�yQ5��`�M���,}�_�"���7�jj��ƛ&���eI$��˫��$��Cjn}xhf�?���� "�`|�D�$�����p�@cn���1�����m�k��+���� �0����rr��ss���'G���t���2��)�L�8�W�Gsz�Md�&98�s_Uv�.��=s�e\��w�������' ��]7_y<��X?��e+~�!�����=`��>Ҕ��s.�����>f�$���Vs3����X�ai =�u$��?MSr��/"Nп�ZD�s Ql\\��1����64{`��k?�!s�͌c7_�B��S�\�<�~EW���"�h�Ty���ћa��$F���%�6`K�FN���;<4Xa��P}Z��1+mvO
�P]?�������E
:_fܠћq�	�����XCh$(��ް�*��X��x�n�к�ty��@��g�=�7��F�~4�I�۲�E�8]���(V*/�,�a�$;~���&_�D��v��ьB��Yû�ES��Ŝo��v����ʦ�j?�r�;kLw���u�fW�+�b5��+{��7�$��R��]����6P��R���\�]��'vH�W*2�ɩL%4=ߟ��2ԩde��ӑcC����n�ב�[��ւ%�S��Q||��H:��֢j� ��nj�(:&?:k��YW�i��A2c�7n~�/���ds�}
�8S�]#�"�{��u?d�!�5��kv�!A��b^D��L6�N�J03ݙ�a��!��?p��p1��(T��k)�U�j�M2���0���VEN���:��s+�j�B�B���U���ab�Dq�v�>���]k���gһ�p(���ޓ�P���)�𓉶6l�{]&�]�x^�B �Ok�����c>��}���Ɵ�u	5b�����}�������Βj�֠�#��a�.�F���E3jU3�u��{e�uM ���#�G[��QE`HIZ�����fܽ� \?�f3s H���#��*(�z8jq�&�i��l ss� 6*c*z��t�L��Rmw|�$�b/13MхgP��	9��P�6 �o|e�^&�@�1BF��1s��Ŝ#�\L��)F����Ϸ��B]�\��y�3�h�~���"���"��dd�YF�+��p"�PL��ά�|� ��#)�n����?�w��f���ѷ�d;�*����1e��$u��lf�6Q����k>G�|���0o���S�m���}:�b��#�zHM�M��)��Q����"�:�R���H�����	}ୁ��0�J��;��9��H�a�:U|���0
k�ݏ�m4���X]�?C�B1�Ḏ��N�m����Ll`�8�ːVvU'�\����V$lU�o��QE���y���>r�b>��(�2=*��k��I,��i��^�r��j�����W�U�I�<��rc����{�����L5�fc�/d�_��t` �(}~L��,q��W��]�0�F�����E_�T)AU�%Ŭ(�(��*���6s��X�y���3�������`A���ؑ'���x#{*���8���z߼�
m�"�s�4�����82r���"�X�-|9"��X�z���c��G��E���%��ӎ:�p
���8����k���5�ibK��"~��M������k���Fv�tw�Ai�ox?y�A�ձ<���h����_�}��5�Ⱥ���cb�Fe<�T�6��}�X�^V�|\X��j�0��M��"r��~<.&���x~b��^�������r���N�"�u9zV9���WL���#��8�w�e����uhk��c��O�2] ���|� ���Ҋ|��"! -'ʀ-2���*@(�A<��қ�A2!�A������������(�K�OXU?r31�-�̜ĦqL�:z�h�NH�W�ࣿ����Z�c�;����희�M_�����vԷtew��ȷ3nGJ����)��dS+H1t�1���[��Q�4@��c�2У�q4s����H�R�v����&5�e���`'�>�0��y}� `�iң�xR�
��.1�6|�`����p?�b���왽DId����ܖkm�&��v�AFX�ڤP]+�>�,�}��?��C�h�-���PHE"�����EU��F�*q]L�n��ޢ���c>l�hd�]���z��zNKG0Ag�&�oAu�=C�q����ٔ����.O�AY$u�L�R�<�'��)H�V]�ԚV���K[K �|Y��G(}��L�Q@ �䏻��2�&�E'�h�<
�$��$?��O\&(����_!l��>d4�bK��KVqji�?��vg��w9EQ�:�#��q���k��m���l�\�Bk����|s[Շ>���Y=W�@	8���+���X��`��؉~��_���$�C{��m-`���za�\��E���T�fk,�9ɣKUս?&��f��H$d|T���̿���p�GG��1��v��*�����'���}������V$!���" [�������k���J�1)��?cYv���=���=�X��ޜo� w�бe�ۙ�	����GD6�5�Q�lu"���@��o��V�	�?^J�.i+��WN/�Pl9v�:kYk7:	��o��ˈhZ���u7i0Հ����(�{k�U�}�o�f�}[ֆ�W�r��U��A���>� ��{���]hu������<�o���?@�f�R4����}Vg��[v Yɒ��~(h(+�X��?X�eJ˙a�<�U�?ٳ�x�=˅��:��K+����T��0� ޹��ժm�e�C����g�[g+��d=;��'�ema��}�	ʋ�G���̇�H�%������ĝÈ���=[�fQ簓t��r��KO�����.2*��mn�H�Ę|JF��j[n� �׏����X����ՙ�y����tld�X��Ƨ���8-+���3[��֏��mE�������\?���W�{�V�q\�g�r9�4���,G�v���j��j�6��Q.��{.n=��Qrkl�}R���_x���RU�D���[����ҋ蕀&��G�?H�.B�(�p�p���X�q
i7��쑱�\��k^�a�ѥC(F�" 2�b�@��v���^��{�c)v0�Г���=�剎�$ś)���_���n�@�Z�Ԃ��&y�B���amN����UE� q̒ Jz��.X$]��̬�y�K�Z�լ���Kf��ז�P�O'���#���jGU�i!� U�ޝ�x|@�L��O
i��&4 ,�̉��r�=`�R�D�F���t�WK�	}�S�y�'>�17w
	�����	HmGm�����ֹ=g�*�w�S��M��y�O�iz�gn�<��=�m�;����ף����>�
k�!��R��Qx�G���-�Lz��!�A��,�r
!���S(�87Y �
��T�!�(b� �$��9��]�0���>���7����o^]�����@$[^N�a<jk(�$9����§#�>D*Ȏ�"��L����F3#G� L�!����]�յڳ5�|���>��t��ڊ����<}8��sjl��!Q�r1�Zz�����k�����Y�J���,Ga�	���
�2j�U����u�]QP���z�r/�Y�$@W��k7[=��'hv�p"2�A,y��v� #POrP��*L:�ʻ5�0��U��@��CÐ�c��Z����o�ֺ�'�~�SXfx[�.�s�)��희�g���� ,K���'���t*�/ ��n�г���}T[�c��ʨ����b�6��w�bw)mq��Uh��\��~:��;q2`�$����0���z[�݉uD��X�V�����1d��R T�� <~Y�d��ĞkH}	A�&�e�Ɓ�щ�N�
ݧ����{��WéZi�s6��{mOL��2V�m�zh${�>X�C+��O�tک`����WW��pt)����)�w�E�f��g`�+�N����nd�1���Q���\�89�O��_������y�H�������t&�c��-���Q�2@���8���t�TP|Pn0� ����Z O�ǫ������d��Яd��VT��ۊ}A�A�%���B脜]1��s����dߎ��X���Rc�,ڲ��������w�5An'U�ĵ�h퇖g6zЌ@��%Qx>�ں_`i�>���3�t�l�~�K��՜
��
|�W��AvqP�3w�B�P�+�98*	�]A�фD�r�%i0= �Lz�8:�UDf�����3���~�E�n���̏]]�����_�3Wڐ�?�Ĕx�^��e�J5Dz3�G�~�߃Q�_��ٚ�C�䪨A�hG���ו��-�%�ɠ�B��+K()��9��t�sm�=!Q�g�$i�@�ٖ$��]�~�E ��1�E-�Pk{��:�/!Ԁ;���,*jƅ'A)D#��E�!}��) ϗ.g�0�5
����I0�)ı�!d�c�8⻞��K�eq�2"���Us���?��
���q�{i��E�%�R�<��
̲k�O��Q*��\8�6��hq�|\a�ߒ����yHq�]��#J�JC�g��[kt	����>�v��kU�K�
�ZK�7�8����5�C$����l�~�|���c����I����(��r"|����d"׃4�����d��*C�y�o�����t�aN�%��7�[p��ߦ:���`d�|ݛO����!k2���W�����ԕ(w����g`��U�t�VI�c�"4�R��=����v^���>�s؟�� D`�|�!z�>��&�R�'�}[�h�6/:ƙP	�=(�S�)������]cA���z�$4[2�d�XAv�Y�^8���a���L>����S���.�^4��.�� b�y%��H�RIjz;j��a6M�^�'O~��&�tE�����;3��g@� DA�A�Ȁ�2��%���-������t|z�Sq�6�8����&���.��Ӝ�.�_S�Ű���E�h]ae�mM�X�T0�*�۝�(V��z^_���E\F�����Qtّ~>�`�4|����^�~�}��Y%��D��Pw�w�=E �Ա�����j���
�,����`�
��V���� ��o��`p@qE�=f��߸�Ww��M��;�� d�s�Q�T�o�z4�Wl/� \��mN�+Q�mdA�KC�d�,'����"���]�u[�[�8����,|��]���\����j9%���v�5J���[�?*.���21"	����.A羋���2PE-��`�Hl�h��1_>�V(���6����Rx�J��$�=(�E.�׼�Lp� *IU�;�MvM��D�*'7���>.G���9k�"��w=����G�_��>�3�s��K4m���o�7�W~���P��4�2�l�J��G�*�V�JZ����R"���|O&/��xq��m�m&HA�'��x�Lw� GH�l�깋�#�e8��a[3I��<&�)���3�K����һ���"#���5�0/����(���ӽ��P��Ê�d�y�`�A��'^=ST���4�qgY�ʮ��_��?��=TرkO�j"ﻯ�N{�rx'0"�a�K�D1GןF��&��gkb�|E7�p�$���p]���F�;x�j�u��J���`�"dׂ`6 �����AY��|���I�jI`�8T�VK낡�׌��L��U��_��9���ll|q�0���i��ht蝞]?�l�cg�^���i���f>`�]n��>b�r�1PC�&R�.�҆��~:!f���9}���x��1��W�r�!)�ЉPk.�>ot�?��1�q+q`2H*ȷ׸�q��\<��<�r�/3��`��%0�4Z͖�ظ�nt�����6�M#J��d�h���xf��v��gS`�9t.�n������Fvǹ+�pz�'�G����Y�w�`�����4b�K�F���
� K��'|�Z��-�a���Sa,A	e;GL#"��%��+���,�����!��#�A�#P`m}�2�-�Z�����ڴ�N4(C�Š?ߦC���?�����:(�ə��N[uX�-�^�L��Vf��V���x/8Rxy��R*T��<t����I�3gR���3Jy��2�"���4�B1��x��>������!���H��B�	��V���w�M4m���(�@�
�f(9�4��ò��G�̎�z{c5@����^qkL7�M^ħ�|��<��/9]�{
B��u��еR��1�����ѫ���rz�
{�N
TM�h��?�=mJ/D��nV�A��4������b�z�/iDlFn��ݮy�/Ci�9豰����ɇB���=g�3�u���u��t��Ӓy��C���t�\:�SŜ��_xg?�S��X�B��n76���r(���-on�*�&�C�L�Q�\Ԑ�ۼұ�ʇ�b�6�'S�-�}�,Gd(F�+O��`]��/XZ���X��]ӹ`����]�)����i�������[��:!2̒���������V�ɝ�(�"�4*�5��q�e�|d�g�Vʜbq�`�B�q.Z��0=h4�����¾���jb�3���pS�dS�g-�/@w[��E�ߕ��᎐�sQ����11"�ȑlurz.�*������'��Sg*�e�6)k��,��bF-9ʪF�åI[��AE�U;6���:�E�P
�$�/P� ^x#ұ���+wK�8$�ǽ=|L��G�,�!q����Z�.���i�t���kD��j'�^1��ƿD�\D��~���σc��N��5����i��A=yU$:��ܲoߗ��j��¢��i��A?v�[�z�$�����cV���K��ݹ�U��o��y6��.�+J�oި����N���_Z��xO����s]�S�C����_K���#7t�
���d�}��2W�1���7�z8*NF�<�w����8Nȉ"$X��:�߃˨n�QS�l�נ�@u @�ރ��z�u��Z8a����7D�W+�H�"+����]��K���Sw���)'qr�,��jY4^B�7KK�����g�>��Ft�ew~��ǹ}3k�.,��C_^4�6=�9�.�ӎS�фa}���U	mʃu�e�S�:�&���񠴦�IT��7L_�io7~j��D�8��w�[�H�����|Ui�?:U�xFj���剧�Y(Ϲ=�������K�i�;��|LP�r/1�=�wpQh�=A�~�w^=-.��I��)��t|��հv��x>V�>X#���u1R�����4?��*��b�� ���7�
��T�K�ZO�q�� �yE�jQD*e-�D ����sKWr)WO3!B:|�8Dq�o��@�6�䉆]���qob&��ǵ�Z2�^�m��)��g_�\�Ш���f��Ҷ�	����
8���ͱv����^!K,��XKg���ޠ\�ڸzlY>�P�<8���/�{2�����#�RG�s�Ҳ�z���;1�$��)q���>��F���Z��S�0���^��銥��\��وA����?�U��QՊ�ݨ��w.�>�n����@3]�M�+��ˋC��r��4,�c�Rˡ��<��ѵ&R�ώ	Mo�<]�ءlZn!�D`�*� '�ұtZ�#��!`�3ڎ)9�a��P����ɍ��Vi�|S�4��k����wHutt����8�mvoh*��%�/]qlZ�v�Z�$���>߃5^�Jl�6��ʧ�4�X�+�w��݇�غ�uu�����G�h��L���Q�;�@[8�����;�t������Px�~Y����T����o��\�8��h�-�� l���
��W�B������!���b)�I�C��\R�W8Ȳ[�ή�CLOn!�%��l;�ʍ��_���o��G\$]W:�`��Y��
�$�����E�i�Ł�oo��E<�8��قR@	f7����zyPZ�@���^������.)��A�?� �Ɩ�w1�Q)U��wp�5E�]���@��G��8՚Mp��ͬO���s�B���Qi>]��A�<�;�aǜ��ݶ���)ɦK̢������T���yEݡt��k��\7z��#�M6��9��*xpm��6�z����D���tN�r'���5���m{)�=��S�*ėh�E�S�~Ma�n�H&+�yŏ4��Q:�J����gu�^#��U��N���\�D�S�@P,�Ds�5�����:��BhB6��Of��|(�[j3 !���m�7��OnH"��];����1�P���J��i
;�^ɧ��19��"�\���b�y۠�_�����<��6��)Z���OR)�[Z�?�pj ���\f'��9�#��<��=臎[W2�%��l��_~[dt�Nzm��|ɑ�C�~��1l^-�m���\17���-� ,���2d@kUXǙ��t��kJMG+2�h�׃��
L�ǃ��2/�X����G��M�"(��.w��D�L$P���W؟����9�����튄u�%�a3��dQS_�B�?��/�Tq��6��.j���NG�n�tٸ�ށR>3�{�Ua��"AX�h`w@*&}$.D���mƦ��RЎƢW�NQ�k�+Uq�
�p��{Y�@%��W��K~���t�D�>�׻���0��m�B61����Ep`w��;N�^�4�+R*�>~)B��8:
��oIQ[���oC@T5$�'�zF��\��&���D�8 -�_x���6x9�*���C��%��=Q�o�����E��m~�o��	������4����С9��a�O���O�ޚ���\$�<�ZY<Y�|�@Elp �&O%���ehSK����I%4:(
��!(SG݈6I��Em]|��j���VX@�b6;iGDD\�G�J/11�Ђ��N&���n�hMq�����M"/�5P��r�Ԍ�T�ٲ-H�����kj䲙��3�8��㝗���jSFUd<���򉜵��N���7�:�:��>�'±?g�<�;l�*hChN �3M� @��}�,?���2����f� �?�=<}��$w12�6x.-��n%�j��]�=��K������'kiN�g�w�՗�7Ӯ����7(��h`�R���i@���a.L|SS]]���%����TW���SSXK�Ԛ���oj`(�䅤���*k7+��M��IH9�ֲoy���}$�f���1�a�uP��(p(D�>�$�	 V���8���ĩ���љ�ػ�#L6z-l���q9��G�N2�:�����9��] .�w��:����$���F��w5d���(YoE�iIX��4X��hN�9d!O��Y��C���1���&5ض/�vUg�,]��5��ևP�]�$5|���#�y*�Q8J*����WXX_�a�K?��F>
��Br�'�	dK�\ⅵ�D�g�o
kk�Q�[�����Џ�Jʵ��Y�31��nQ�#
�?b�P��~�D��Mr(l��~��ҁ���tۜ�X�+�]�J+��r����P�֋���n��&��T��w�I\InQ)=�YS�������v5Z��樃��T%ӜF�P��Y}h�@E���\�͖��@����P� � �cP�t�O���.=�*vT���;�IϦ�K}�2��V �<HpTz�"���w>Z䴜n[�ukx*��;S䶾l��2N�kxo�v�4�¸�}ļA�8��z\�vJ\r�Z��[뱇�I!�f�[-�X�oAh���s��23C�� �2ڞQh�$�2� �1Z���Jﻪ�5C��H��	n.C[��m��9�{ ֟���'�27>$h`�SFi..Ȃ\�"w^"���Į�-׿���������qV/� 
���~oA�C7�a��T��K���4k�����[�v�{	����N��5~1�&��QWx��
�k�TĬ2�A��V��������}�0w�X�o[|b�8(s��C�D�jnV܇����Z*i���R��ґ��O2� ��#Y��|��ot��vɊ�9*鲦{W�ؖ�݈���ғ;��ۥ���,�����JZ0'g]b�F%�qoiÛ�!�;��A�Kֶ����4�<
iM� ?��'R�&��3�O��Z�J����Shf'7�jVja�4�1���]z�ז,���^߄�ѧ&�<u��(�ު
`M���"��)�۝Y���܊ϥ�<v�k ��) �Ȅ�R"�E��c��z�X^���K�&d���
�6�"����ݡ�?lW���[�8ZL_�-h�N8ZkRnx�<H����������>���+JL^r�2�_�L����_,������L�H��2��g!At3�P��d�(ث�xx��)�X�tle�}#Y�·!ϰ�A���^�Uř��*��,z!��_�t�-~�#�nB�x�;9҄��H����׍����nnd�:�-X>]z@h(�H�n� C�V�V=�n;�H��f�4��ޯr$&F6�ig[�l0B����Q�S�ki��S-�Qq^��E��u��0ׄ�Yi���4�$9=Z|LH�3I~q�u�pqg�`4}�*=��x�/��bb>u
�_w��ζ*р׀e�aa�Ju�4��ҵ����-w�
Q1LV���kJ��JR�4�Q-��Ɛ\��{{�g����V�%K%ӂC�C��������묞6�+��?b�q=��`?E��Q��3ţ�k�]���,�o�g�������^I�����s+����Kzf��7�,'�bb�WԜ��j��-�;CɁ�?PK�qݰ��z.�:�����i�ޕ��s]x4tkQD/g`�>�7���_2�����e[�`��o�!l�Ȟ��2���sa�C	��v�l���mI��֧+l���yh'�y���70;�P�^Z�3W�`�0��*�� �U�?�w�`�H3�Nܚ@�]����@\D\nl*��N�u�*ͪHܪص" ��5lF��	���#�����.J2JF��H ����z�'w'�5���gI>�Hvv�J�;��P����A�T�U�6���lGf
i	7`wIT�29%����#�t����і�[�Cb��sօb�"�W�^ǳ�y66..b��Ӷ�	����M<�	)�֬u�i�n
e��2oa�B��H��V�Axw�j�����3����u�U��D r:Ι����M�ˮD�t����	�|���Db�����&�L�gRp  }x�a�8xx�z]�e�]^l���ѸM��BB6�3:�C�ǳ����)���d������zU��e�X���<zҢ�K	w���FPϺo!�{#<�(����7W�W�Q��W-W���[nd�u���/�*b�\�e� ����~g��l���ޘ�����?8 ���+�m�q�iz?P�i�yɽ�������u����Ov���_|3OT�B�@ �W\�f�}X�y\�B�t��LE��wWD4|��~�iq-� {ZYk]��>���]�䣧������0� �R�����2A3�qe+�e�g8�ns�/����b��	�����)��$����a���?5���f�k�j@�-ŕ��gd�2��.� ������F��"���=Z�ˢ�} 91n}˅b���j�@�\=p��Ԓ(0H�����V�rփ�?- ���Y::��bb.
�*���~���R��5M����k�kWR�,[��Y�~�~�rE�{v�rq�ruW��|���BGWm����� �E��8y~�}\��_D=��0H�a���^�ƍ��c]��C
�0���m/�7���of. �L\g�U���R���2�;��u#������k���#�� I��m�ٽ��Պ������!��kb���ǅ#P����Rꬷ<�s�w`PTYC��UfY����Wu�ܫ�Ĳ")��$�܀�Z����0��Z���o�`��q�ܟ�2�b�z=J�qƣ(�Z�՗B$�c�6ȣ�㳝0_�q������:�����3`��e_/��j��;#�����4��?�)��!�W��鏨	C�0 �4�U�,��#8⭯�](xƵ?���"6Z��/���_��U5 GyU��>F,��Hsb\�E� �D�;���(^k7+%>\�	
���يӋ�ɿ�����	��{oA�����e���;�"����/f
e��:d%�l'����Gĝ�q��ft��j��Y��g�(��;�	V�pG6�3یE�ǃ��]y<���`E��vX)F	�-��W>��b��xJ�,�uP�q��6H1UO�UC<��GS�5��$!G����\��1�Of8���:�3�JMxU\Ƭ��[��|&J��"ô�q�۷���	*�쭨 �BV��P�WFZ�lҔ9�0{�d4���>�J�����0���/��{ ��H��)�T����9\tWi>�$��O����.D�b��̉|i��(|o�.ԕ�!ޑ���~�.c)�F��ݩ^=�S������u���YB`�����^�q��*]7ɓ�O�>�+ǖ��S�iN�^_Jp��x��,����_KF�y���/{;=��:3��9BMv���af�^�d �0C�i����	�5��������(�gЙ�y�X���>o�6<�d�:<����ػzC����Ć�:Z�(�n��e3�ҟ�8�_�`�Px�u�^��癘:��`�1h�
���fNZNr�#���8O��ҧ�q��0��=h�7c�����h~����ß���$��yv�P�_�k�������x�_�X�ڮ��{�[ؼ�iҰ�~3M��~+熮����9t4�y��>(L8�@�Bfc��>.&t蛬�D'NJ��E�(��'�g�� �M�%�����x|8̓��=8�f��,j�y4�j�ѷ�$�V7�g��߅��>�~����l��)>D1_�>�PR)�"�����nᛙp6U�m���hu/1�m��?U�߳?
��3���[5��ip�Sط��4��vq��@XΘ�C����K���F#]*��Q���4���"��Y���� p_@�b-��3L�)�h�>�����yũQR������.�D�*�v��D;�I�gR��wہ|����6b��YS������v/��Լ�����7R�0pM�+���18ǰ����4��E����ޏP{{0����g�Pj*�^u%�dKU����&M~�Q3�ad?_<(�AM�p�XǮN[����4����c��3�+I��
`�L�Ď�w�iu�԰�-�,R`��m�_��ڛ����UƝ�@�� )�5)�s�ק�T�@��\
't���p�OOs����DVb2�wn�����X�Ǖ�fg��J������?��un���÷�5q��u�*��V{9�*��S�N�=�9T��
k������{��F�kc!�Ĩi��/W�ŧ"�Ůw�ZZ��ƺb8&[�ה��C�c*7Sp۸�{`&�4s��p3����7籠������j�<�������̀l���1#��F�@�<��IƘ��0�`�'Fi�e�/G�H U�w_�uQ�4xY�裍���1ŏ�~nk~����Z0�:�{m��|[���F�|������M�]��ɮ{�H�~��+I��ҟ������$�JB�˵�ӟ��WT��^����^��LRg��>s�� >��6=@_�>�����ڑ��� 7��Y~�ȷe˥7�7?�����Ae�
�d��x^��I������݈�8�*����گ`���	��BBl�b0�|�zq^�!�������a�P��D{C[�Q����j�D��R�M�q�����v^�3��O�����2�LTڙ�9m��8�KW���=���ne�u���qt���w;��N�ivݵ��ӑx��-Ɗ�PZ�Ž�F](Q�7+*��O5��ݒ!p�=�D/��4���0&ٹ�{�n�n�Z������뭣��M�o�o�����2�jX
�I��z2%�_���*N������n`�=p��F�kNǜ0_�ϐ:_ۚh�u���<[b]~~Z���mJ�G�(HV&�_w�U�V�%�F���c(~�����7cWb�nZ�s7����<��H���5F �='�=�Ikr&�@�V�3�����@N��Z�w9��W���:l���"�84T�޺��,�vWus�-�|�{�D, y(<�uޛJ�e�p;/������Y����Xd-�M�W�u5AqtGD�c����W�l�8���'/ւ�uۯkgErd�|������.�r���ajM�Q2eAԶ�\��׼}�æ&il�����i�d�x1^�5ka~�\o�)���[{;���d�����K{��F�NC��$�q��3�̇b�{J��'	�7@�s(��u��]r֞��b�u|��{m�
��Q����\V��7"��p">�q�&r�,�����RX>�Jl ֶ�u^���]AZ��@~�����>���_��������FS�7�!��ܲ>��<��Z;CC)A<�I��i,���H�ӫ5���y��\�汸��~/ր��(}b���]��lF�&�����~/-�0�y��E0��"�p�5�����+u^�ꀲ7�SyE�~E^���N�ȝ�s�o�`��߾���$~�V�[v�y����#��ध6�Dץ��3��!׼>*d:�������K�.,n�!������L8�����SEv<"��Rb��kbE�f6�o��%��膂�6sj����1{y�$ٹ�=4Ŝ\"+س�	Wk9v�p[��-����jxah_�5���&��͜a͓�O�����c�OZ����M1c����Z���g�jh�4 r���BZDU��J>1D��ԌHҁ�P���jg�Q�[���l��	p��TR���z�>&�+�cF�ٯ#���F��q��l_ܺh�t��l�Z5Jk�.Ԯ�Gk��+V'5J�M�-5"$��{�bjě�_��������=���9�|��{q�}�$�&��nͷ��т��=�_�����ce�>�SR��MV������f�ފ�VX;����3JH���Y����\���o[3�+_I���gnK�৩�q����+ؾ[��S"���j���l��j���"�@����?]6�h��3��]^R�3�E �]�x{���+�4�*���1��(�Tb7D�l�E�E��D�`T�=Yk�f���d�˯X��kn1UV��UԫX�5�f��D���!�EU�$�$�fe�Ax�\�;��A�R��T���h�1�qΔkn��|��R8��n-��m�pP0��y�	��}���D����s����	F~�҇h5tŞQU�Lz�?݇��������F�&��Ov+���~�e�EdjF3����8�跎��'�����*�/�ԡC�
,��|H�D�3�I�>
h����Q��.�(/vC`~�������_�0^��e`p���c�^�I�$s$
�a�s�$!y�3�2�G��{qsL���TZ����V��ҽj i`��ь-��6/LM�vؼv#�MO��8*2���	������U���;t��nF/�ͭࡌ���E���G�7������+T�-��C��/�TW��^�uѱRs@��=̇_��]m��E�R���U���|"�l��f��ڟ���TF���~G�n@T�+�dХq��~G�_��EP��j���_��&@]�Ƚ�_|�b�^��N�?���'c�V��ѯ9"�[�Pn�'�s$���'�p�-�,��°Ê��3�5�~�،�C��\��VX��?�X��s�bw���x���X�2z�%�y	��ڇ��%D[��#�'�V�X�_n�?�r�ӧA'���OE�z���̙�;ґ�ג����|`>ĹJUej�'����k3VeϮ,�,�����47��u��O���p{}n}t	�������RD��y��qN�#!y �ƚ��~����/��`����i���k�3���u]�_h@��2;G�ٍ]C��_��E	b�~��?~O.D����8U��X�C'��}�-����M=,"A���������&���h�^ǜ!i�;��I0Ƈ��h���O��g�/�MH:�q��=���qg$xP����?�m��Lz�2��%��e��v�J�E|��D���g�|Л�W�c4�OuA���3P XAP��$��ր?V����^��oXި����-�gi��"4r��SG�|Rx���S���}ʈ'>���S��P�/2��#�A����E�����||��?|)�K��,�V��f�F,(#��v"�S߼FS�d�EI��vvv�J'��'{, 0�Ψ��RX�,���=�/8ˉK��\!!���"�'a�\����&��s��&h@�������X!#wI�.C"�-�JNIQ�2�g��s��Ntשּ��TSoF�XѤ��`8����������k_�f�>S � ��e��_SKI�2�Arn'Mo��KI3w��.F�L��5��9��mӉ�|EH�[��#��L��Y#�Ѕ}+2�R]O� �fE�at�Hyk��?��'������&���Ɓ�E:�y�T��k�4�T*����-&��^x�G6w������c���|�F�۞;���ӳ�/A�Q1	�HOt��f^%b�h:b��ԋ��PVsPe){r�ρ�9d�S��XW��މ�7��}S�k`X�ɫh��U����7
h����g���T���^oڙ�Y���:���[�p�L�@��㡞��W;W]pA!�A��}�x� Ʈ�7S}}��MXw�Ӡt����zծ�鉏����|̮��IJ6��4cvz@3���(oq~g���.C�1+�������+U�n,�W��JU�'/��l�������
 �HU}��'sE�~#u��z����k�oL3�r���q��O|�uE�$S�юb�_���Ӎ��Z&�>�"|���1���yXF�\N܂K%�ޭ�ٜ�L���吵�ک�G��@�]�a6>"^
f�P��8Ȏ	�؋�sB[%��Q2輡���n�W�^�Oݤ���pmn�N�k���Q[ݔ��I��M�^��&���#%�;E��v�F�똔�2|�QJ�K��'�ٜuڣ��M�Ճ7��u0�T����\�H��';x��^M"�v>� �.�G�������}��H��&�}�50��n�����NS�h�B��o�`R��7�̰�0Ϳ��)M�&7�����i��_�'-}�j�б���SD}���|�bZ���x/TMP�7>�����4�6d~�<���;��bP����$�y�K;#�����!Щר�����{�S�H��ɔ��lt5b�|x��'���UBĂ���({�ͥ��Q��U�����$d��L��2��cό�$���~W��p-�֋-*~譓 	Ik?�!Ľ#�~��E�%�W1�G�N�w+��Vj�9��'��Ǣ���\3� 1 4��k���k��Xv�"n�p	��k����7{_����~��a�t�*��rHc70��*�p[�/�w.���0�݉���]d�����np���k����/��~�[w�!�Y�v�J�BܨƫM�ؐ���E���� en'�d<W	1
��e%�!�s��ԈG�G�>����?2k/�$�Q����K���:���y��6l@�:MUiͭ�1�� ��%�� ��a�n�j/�%����0��S#�����?M--��,|\��e�6���w�2�Ւ�.�Yxp|�����16�{p���O��Ĳ4d��Ty\:�uO��)}�X��$���@{˲����	���>sc��@�#�&��[v2u��j�ٶ���Sjm�^��g=�V r$��x-�5�`����UM/��.�{�Z#٦2OOvڥe�l���v�L�2�����W�[U��v�����Ҁ��2!	���z���R�4]�����t�^i����
&�Ԛ���s�̟�,ĳ(��'�~e"Y���/dC��lb��W(��8,���!��WU\nj�9ܞ���bP��fH>��ڷ�3�9�I�+�	ó͟__���p�cz���c`DNj���e U��F�Ү����I�+�'�2��/ �E��Uv^?F�U�E�}_d��⁪mt9R�C�`�a����od1�l�p%��
#����zЧ�O���h&)UuOy���bt���=s�Q4y� ���,�D:�44�Ш��qħ��&�ʌ���aא���+�c�Q�}�M5k�ku���2�����3������÷������Jʃ��u����.���;�W�}����I���U��ҍ�
0u�`_J7���_Z!	�� ��_��	��(.������H%j�%P�Ւx��A1�b�CԒ�5"[--�-��'H0-$"D��x�K=s�FO;jv+��jy�����ϟ��ɬ�f� �M侯 �����\Ԃ���	˾�a#Z���g�Q��B������H��
Iz���w��kt��J��޿vl�c�&a�p>�*��B3RDMѫ��.�,��_�!	.��@�P�����z~�K�����X-+��l���Q�q�vK�D��
Ƀoz��b��nŪŶ���,�2|Z�m|�CLl�K�L�������J�D_`�Do*ДhQ#\d'�z�b�"���ǴK�f�;���:����g����}F��\- +�l�O���M2�]�sS^�W�V`J=Y�Q�Q�Q�QG\�u��7:;o�dw��C�L{��`��h��K��&�����K��/���<��?�@"��_I��d��?
C���x�. �Z�ˇ�J����s��9@�K�{�F%?Dy 3��}������%�� ��E���گ?�?O�l{���<-�$�!�����C�D��OM���'

&��<���s�)2��˚A�gß�K�r�$X�7�4)�Ҳ5���QȉZ6hu�J����ؘ�ZW>A��%����렲D�<ekb/~�q���k +�%�_�)�*�U���2>C�8�(n_kg�s�LԲ�A]�:�%�M���ք�����ܲ�8s�`��$ދ�����cP��;<:��I,����9	))s�g�	|#��������PXZZ��_�Qy;u�����"����m����n/�.&�E$Y���D� `�ѹv�;�I�Q����kN)}��3%��w�T��]}�"�k���}�T��6�x�y�ϗ"#��G�bt�Jd���o�~�-���� �a�<H�^�Ѫ���o�L�����Η^ �����st�#�nSni�?��C��6���y��9 �Q��Ժ�A�r�y�����s������i�{=�=﷈�:5�գE{d���H��#�QЏ-���O�{?S�rk���ٍ�1k�J���cEo ���H:���9��bi` leOD����lH~�a����mq�3d�� ~eڪ'5������)m��<���nx�f� )���#'���kP��\Pm;�9�m�o�沋�u'W��k��I�Zw7�"�-ն�8$VGA���C��'v�w�vU��g=}@��*�Aui�[s[
����(������"�7Z�,j��س����jZ��.v%��$ӗJn��4�����Q#iꖜY���?���;���'��{��b�d��d胣�m 9ס[꾏sbѮ8M:��y�5R~u��x^CnE��Μ����*׮�o�%���UD��)\:��Ȥˈ���Ӧ�n��۔Z����=Ǯr#"�Cvw;R�/Iu�, Cm�������Dab+�8�,�ͻLp��?vI9>4Fr��#֊��Rm����Ɋ�53�ĨA�6���\��k�r(��^�+v

z���A 8;�Ae�ex��ϳ0����|[��(��⻰�*����"���m��<��R#H���%.�2A
 �"r@�.��R�M_�}�Q�����|�(����_ n,H՚*
�[y,DE-��Qڹ��yH]x�W�|7��o�G"��������K�W�@[%����z���~��e�lW���L���c2���\��Z�O֤ ��J"�ӿ�����Y����@g ��-(ic����y'�T�F�*u�_0�#��, �P��_��y�Ň�s#:�OM�j��Rej�uX�*.�>����=���~_���c` Y����c>��U*d����_��\S3��xR�Љl�?2Bih<�h�vL@�S��ҫ�~�N{=������Ut|�g��
�yW��$53�6�oS{Z��/cuw�Z���{]]��Ȑ��M��_��N'��?*5hԗ0Ж����WD��G��C+����-��.�QS?�+���2������SA��l�Txeq!��V�h�0OK'��:��PX(�7�a$gc�mV�5�i�-�� �Gd��"��p��uO8d�x�5���#�$x��3e�:��ݬD��Y�8���)1��O�y,Q/��$�����Z�:�Ěo��X����#Oy��8�Q�c<������7y�J:�{���I*��|ퟵ�5׍k��sJ�֖�G���������O���;��8��mcl�n0R_�%�Rq�S�v�J�
�����}�?���I��U�W� ��]A����]~<�!L������+��'���cMnC @��޻���[����5Z�1���+��,S�݁�Ha�~B��O�;<'�b����F��{c����ˇ��o��[+(K��w�'/�'�!�5�з)�R��	G�ݖ�Y�C�tUϩ������C���Y>ͫi_�_�]Mqh�(�2��k�����`&���Z߻�n��A�U�!o*���R=������%B	�vc��q4�i/���'2�Fuj���lV/J�}V#~��t=[�ǫ�I�[U:d{����l#>4���I�/�TC1We�2��5;'������`��r��hf-�wˡ^]}�x���oipA�ƚ�y��^<m�Nc�J��Z�CyE��9���6��B�� ��V��C��@����	�x��_�J�~+^&J �o�I������!{}����B^&� ��m�`��(�4�*���?�2�~=I��/�����H�6��`����{�$�����-|���.4ԝ��Kڼ`TBL�:��q���E�{;ŋ��	�����jbӥlmlt}��Y迶̻@��"N��6jL�u>�^���H�22�GG~K���>��� n�N�u�Sw�82�IѦk�Q@�;�"vpi��zc>4D��}K�O��O�ͷ��^S��Hy��m��U��Š� ��]d=R}	#,� t��lEIY����%c,���?NO�>�)I̻&	��5Y�ɭB 
�`�p�@�θ(��v7�rRSj�R̕;������p��Q�?�rw�����{�oU�4��"n����zmr�����'��"I�dޓ����/1;�BE���4�dCL��E�#���[�,���`84�c�(�׷'�E�[�����e�'�J�h}��Jz,�-S��AǛ�$�E����S}��6��0hd�C"�ۘO*w��^�H�b�������E�E���ݢr��Q�Rw�rD��)�CV�o��7���>l��j�S$ڛ�^�U�%nʼ7�q�S@�~���O�7ܤ[6C���	ȉ]�ǯΊ{,a��D�M��Ř���[�i�si�pӵ���K�"5��M&!�ĹAK@��y?n-,���D�0�ɷ����)k#h��?3YO���fg����<p���ܷ�.40�2|E7�I��A!PȰ����|z?�'��{	���(��'�����,�|Myϓ�KWq�f�����F����qG��=P6$���o��A;U���	ʪ�W��wI�VW�e
 Wg?�qPV��n�p���\L{�P^���Ը�H���a1R��"i�
�'`Y�u�xpO���*�go���{�Gy�Հ�)R�ē�]�:�9tg/�ڧC�xq���p�K3R1����L�+ݳK����t��=�
oɼ��+��4sL˽���{}-���WH���<�Ʀ~��..�(����J��H�>��������dk�F�
���<v�>�o�����{���B��M�0!��uX�R�Ǌ|�>ߞ�T��̖fLD\�������ϩս�u����~8��mk,�8�ya~��"Z�5���N��Ҥ��Ur+R|�؆��������1)����	Vh�75jq��=̃���|�iOy��A����ӡ�7�����5�e�곧LM̖�#��y	A��	V�f���Ve���m�����q
�.D��J�^y�Z�Dwnq��*�q��'j�Z_UCNv{e~."����ռ�)ڱ�q���E����H���� ��4�*L���T�}/���]4����R̡��rӌ��e(籏�ܦPk<�]��"��ne.9��0�U�o��������J���[��ԟL��ѷ��1:.��L���V�g<�� ���.i#�N#��-�����I���R�L�HGF�����48>��.���:$����Vm$rܫ��Fi��ōZ���o��|��̭��
�U���T����+B&����}v0�F��Կ���a�`����М����J����Zϱ;��~Ǉ���`���Od{�I��� ��@N@hV���T�����4�?��Uh��U��qXw��9 �E>1����+���"LP�'��qpS|�^����0�h�o !]_�������QH�	o�< �P!5rrT����x�Ń����#t盏�[���Wg��"�#����p�� si��"O�cK	�g
L��^R�����Ga+�b�nG�A���ʰ�+��� ��Mc.?L%(�1G�!�m��N_P��Ф�1jv;AtxnxP��9bH��?V!<CJ�b��\���O.��/�UY�i����s�L[��V��;6�xR�����	oD��GE�%R��%��-ʤ*�0������)�jđ4��DJ0�����|�.=6�o�X������n���8>�8��������4�gR�<��v>�b��xV3�]�N\hx���tT�Y8[�h�84�B�Z��N��c��z�R2Vro�6�o�ۨ���NnC4p�˶<����I��*@_�<�N\K!t��t����3Y_�h�K�b�����v�XD��3�HK�?��_$�b���4cK:6�i�je�8��W �\��+f;���9�{�²h���w������R�z����վ��7m	mpQ���\�R��Ɣ�Q�@_��7��N�n�F}��m*@���j�Ԛ�[���Y.�(tN���Vn�y�R'3Y �TU	X�G �j�*�yÙ�K (X�Y!�C%>�D�A�џ���>U���]�6�϶mF?�)/�U�6��̨��Tſ�ys��vx<��W�t��!��Ϙ���N�w3��	�7��Y��V��]�SfG[ۆ=�pj�m�K`��r�����N����XOf]��[8)�����u��o�]-t?[��4x�n�~nƪ��l���`�@Z֘^�����z\½�n32פFv�����1���W��Y_��'bL�H�se�$��'�&y�7�t���S�,	0�Cn}�����a�w;$=.ب��g=��UD�H����2��*-�I��������"xk�	p��n�X����3�t�[��7��u%.@;'�X9	3f3ϸV��czd����2M�~E*��I>/���`��%S��֡%'��"�T�o�,=���I{�km��E��O�S2g��z&%k��*�cU�T<���K'2�j@���� ٿ^�!*-&�F���2�~
�[J�kT������Ҹ��9�u����@��i;�Ar���G����L�徲�'K��r�xm� ����w�9���j�������͝���-��%'�yg;A6�.��[F)�����{%�%�����Mӓ|]�c1��a�)��]��T	�s'Ӏ�(�Ryo�ı�ʽAi`�"��{/��K|1�rur�QYQ�}P����x#��wq���~{���2h�U;��w�� �8��Z��<�ו �4}@�sv�:���G��U���r�~�v���~�MX�>d7I��r���EI�ܜM�0��zJ�Mޔ��05&��%1�����82Qx�?�Y]�|�dk�2"��"���n�=��j� �;��9�@����(*��@��L������B�87�����S_��G~�ǫ�� $b�EZ�c�n�9)A㋔@;�,o����2�9�9��u��C����Y�`��]Ob����H?����������r {(�r`��7n����Zm�&	R;�)�wRRT�a��t(B��x������[2c��I�\CB�<�����sf�˘H|��g�֭��c�������<�b[�"Չ�֜�HY7 �w0��`Rt����� N��{�5$ �K��Ƃ����|	|�ƅ	�J	i&O��	�܄DF���r�Z2E��լ�ϾO?�I�����d���v{^�f>Z�a;��+;%�*	̓�p��B��%yct�R���y��L�q"~�-.S��Њ]*��V����/�<b�����?�֩�o�?��V���A�����=c��ܯM��:�C�?"��w�!zn�^��a��B��۱�x⇮�3 ���k��E+�3�ֆ;͋�7ed�=��D�{�\����ŵ��:��] �Eo]�����'&�J��/Op��@V�$���li1a�E�(AK���j��W!�N���Z�rV-��` \��I������E_�z�g���i�,���?��1�8�w�qw�K�0SH��7�����`F�K���,>&S���YWؕ����LeE�_�}���D�FyZ��UҋV��:y.�]G|�Mŗ���7R�݃ ���rV��ۘ��Lg��ju�L�Ru�;ӑ�����-��⁲��[A'�r𓢆�@�wNv���*�
^N�%�� ǑG�����23��=�bC;�)�	w�1�8O��v��`�	>׉�s��mZ쉙��b%����*�dm{;��g'�s�C0��'o�@$`�Tfu��0Ow����} A5bX%�]��eW��汨һ��"a����=�v���%�N���$y7n;�QݰwY�¢	_/)5)`��3愁ЈE�ɪ�C𛻽L' ���;nK'�����·�j8���[�)�c��ǥ�S��=~`1g˚��=?��=��<Ļ��n�'DZ�!a��-�]L�޸`�-%L��Fr��Q�c�U����h�G�*f�a����驰�k�S%%	�;�`�2�D��P�V��"��GST{��\N^��{P����gN9}_ii.���;���^�^���맜�j�U!!U#+L�6�V�ţ������?_��y0,���#p ���t��@,���s�F70�Lg)�x/)Ö��i���M�_���ŏ����]�	�ʫ��3���h��(&n�����
�!Nr�b6m����_��p�#j��c�m����-�N�O\x[�ӵr'�;Ղ*��"E��_*k޺A�G'�"'k�ɭ�m-U>t�swmt�'@X�x�TՖ��&gw*7�;��z�F��T�;��ѴN5�o�u��]�Th%�U&���ȾEB"*<��d�NwnH�jq�5��\�}���m����?���Y"ݔ6<|����`Ny�{s�0�������j�2f `�t�l�l�w ]u�͓��Q�� P�o4g�O�Kዌ	�����'��ï �g��.O�o%YyR*�K�R��{i�:��[;� 5 �QYH����rB xKTjX��(C�߲,�e�k?u��{ӹ��!tr�=�pg-~7��}�;N����p7z���%Uy�<qE���b&.$��^F�c$_F��hwN\��%Q&��S5��-����	�E��]a.��3�Wr�8)�/W9A��f9����׀�.(,a���^O��[�gӆ�j������ڠ��pǒB�]��x��7!�m=Z�]�w���'-W*t�OJ�S���nU�ޟ���qq�d_B>mJ��[�8�-|�����m��#��/����N�"r ��N;,�wr��g^�ս�,��DS���Nfk�Q��5ٿ���۾�� 0�i4�f^��%!�C훡E�Y���ϧW91<�R�V����Z�M���=�e��Z���Af�G��+�K�\�
�&���|
�L5���|l<��'���u�R��R#�H�jla��{e����p���=�C��B-E������<[,%)����[��R��m�B1����YC�9�W�����QlWQ���v=O"pPkķ��$v:;��E�O�{?�* �8z�����U��?�I79��"<�[ˤ#�L��c:Y�d�&��(����:>��/�w���#�nĪr���eP��E����	S��WK�����49[�#y4�&� "�4b�����t�m������1�C����g����8�+��b���1S��N6,���B_��<P%#��]�W�g%���ڙ���a����l�l��>�ky�%Oh�q�٩K��@�&����/�Q�=���#��]����,$�9Y���L�C��������}�~^��'�x��$k�����!�&�=◈�'��Q����ڵ�Q��\֣�l�W��aʢs�@FE����S���Ă��߄`ch^l`h��wH���ƣ���P4\k0�F��$� ۟9�iU����*�(��66ή��!0�+�!������0���<�ߺ�~*�L��d��
l���̓��'r�kܺ0�o]Z޺�}$�#?~x�G[��Z��OO��n�0�q�]��& F`W��]�ؚI6�X���e�S������՝М~����Υ;G�T��"�[+�U�(P;�!�~D5$���N���?��DP����}s��W�qmoƈ�u�FJӭC�;x�j���f�O�?��zΚ�쾞^_�>EuY�/�o�v%~��[��ڱSܳ�����ط�yo�ߖg��1�D��\��	�&5�Lb�bnڣI`޵�~��}a)�?��$R1zqa�V�c���vA�p���Ӛ�� &���_-�)�`ms�5dSY�"�����4����H��}"�O�-gs�f���Ƽޫ?uM޳<!b���� /*�'�l��e0A6%��X��5A��� )�<�?��t�א@����bZcͩ�$�s�=�I���#��Ӗ�AL5��n��5�0B
)i����N�X������o�c|���)$sA��P]�]��-�y�	��zh��}3�ɬɸXz���P�n��+���Q��z��J�v/��|�y�h�� l�"0~ų�ǻ�6�+�uOg��tV׈\k8�����v����7��D.0�Aw���cz�H6��j�$<�-���Yb�2�ϗ-h�9��E��û�y���ܺ��]Є#X0�<�5I�Cf5Nf� ДX���%�����#Zv��KEe��K�]Wz\�][�X$o��.$b旖�����{d���Kv�!���{�v�$*mK՗��ݙ�=Z'D-K6
6��\Xh���W�a�nm;��w���#1���8���~�ט%�O�u.f5Q&��M��e��j���;DIR��f�,9-7?/�[4t��m��.�pM`�	j�묋�%��~n�i�)�6�ʕ�}CCg~x�	��w�5��)nL��Y��M�m�t������A�p8\Z�e��vv�MLդ���F����F|1O�.��)�9lP���G��{���v�/�}b�����&N���vd������h�An��}nb�G���� E��W����_��EVi&��ֻ����]�rq��߈�����MA���}J�9ʭ�l��\��
-s.-�W�c��G_a�E<�3�&ydG��mf�亃�$�uQg`�K�^pĞ�{��{u�
Y�y[{���D�KW���	���|K�+���2ׇ|i�A�R�AwTj��[�i`������Y���C���zʅ@k)^(O��H|{�%w��K$K��G��J_�\(�vd�e��1)yⵕ�5�1�H.�;�ŀ���ʭK��D��"�uw�f��E3�Y��鈕"+[ޑ�[��o�=�u�$�x����,�zK�Y���X�����*�x��|��l�P�XO�бt!l�Z�P�yL��i�(?��s�C�n�j.z�1�7~��SB�&�	�?���aK��ϋ�q �6>�ԅ���`��D4�Y��W��8~��xa�z~fSZ��DFo�m��4A9�:�����������{C5j��#�ڀG��	)Uy��$��I�����Ώv�}fݓ��s|���mkWk�OTx�gK]��A�tn&J�p���S��F�ğ�`��a����.tZ
�{&�x����,��$���2t�E�m�y�|��"���o����pU��9��ض;���;��خ���:���:`��'�����:3k?
D nk��1]�8���NW��~k��J�Uh����Gm�U�������i�5ҧ�13�D���QmC�鎮D��Z���ur	byr���%)�R\J�b[-�����K$DJ�^���
��d��⤚?"���5r�����A�69N!$j�c��?�8��ٳ���ZƠ��)Z+����ഺ����0�����L��hL�X��XU��V����\W�!C*4�����2��8x�*y�Fo��:ߧ�!�	�ok��G%�;wE&��/6wCv�4�;:V*O3�w�n���憷Q���/��v�� ��h��!�� �x^�m�1?=�2�фa�QX�"򎦂��7ӸG!m�
��a���
�f�%Rg��T����7^߽�N�;Q��>
�/{�܉9ohz+g�����-�]\A����3/�|��3q�G��Xoڅ�������`�7O��b��U��o'ɻ������4߲�q��!T���A5����Z���cD�S4n�s.��~ҧ��@O>� ��=*)!�P

�0��ݯi��_�y�~�2�T�%�Mj��i͂�Ԃ�7?���h��!�Ph�(�Б#��~�VL��\�c}	��;�2�7$ST�!{&�[sy\#�#��ߥ%�U3���K�Ӑ�o�+5��y�H�0m����YA~"B14d՝4�=n���O���ѝ��2��4&�C 9��y�_���6�ӑ�
�Y�暬Q�S +�ǐ��q��ĕ�ǍX;���dNe���w���I�5�KP5�~|||�+��U� %li���أ�v �h���mS�a��c�Sr�pCq�u;y�_�P�!���B@ӥ�1`fi���ေ%�m��?�*J��w��_zL���0k�E\���Vޱ�N�.��Ľ���JH�ay��-��Oo�����QX=�?P�ӝ+5 )bF�^GO�ɗ
�eK����\���+��D����گ�)�P����
�)�z!ϩ,uO�liG���{6�vR7��"$l��9V{�[ּa�d}�SS�%cvx�vu��c���R
��c�g�U���1��>��J���n̶pss��IH��,�'�X�{��4A�
��1�^�v/��~��`�LnS������sG�\�l�>[��6�Z[u��*5�\����8fw���4��Q�S�7��ƣgYe�'���]QX��@P�Q��gs�R!k�N�&~��;���ވ2����N�<*l}|���d�6�H�����Lnĉ���6�/S�GQ�=b������B]{io<���4�HQ�Cq;����%�lx�7f�6�HG���<Z�3Z>g����&Os/b�'@)L���wR��Ў�ci�YZ��qX|�N���Z��x�Qm�}�C�$QZSl6�cX��L��,uL�"�4�w���yb>�m/շֱt8 D-�o�^��!�{ �� ��"�N�PQT�Cn�
H�kmi������')�p����c��7t��~T�-��S�_rhV&��*�{�;�w�\&ZP��W�E���������9���n�}<�80�9yE��&�����c��kNq5l�?�3�wݸ�~��RD�����A�ȫ�a�B.�<)����0"��Aà���E��!$T��6\G����[cc��wW�E�Q��עęlC5��I�r�g3{��&����=���1�:�㌜� ����Ŕv{	�	��ϭ�1��J�m�yt����G�f������t�(z1\����Y>��)G
q�vPWj.4��劰���t|�{�SJ�k��19Y�Y(�M�+񄧜��n�y�R����8h,y9���_�~��[�$�t:1@��kş�/��Ͻp#��:M�����#E��T�	��W��1S�f^��>D?���-�i3Y	������:ׂݦ�MH�d�^��auh�*��f]+��6����_+���_:��2�;���?�S��k>y�cbq�6�����j�bP��Vs����qgT#��H� Ф��oǘ)`��p����������y�UH$�)~I�����	Wi}(V8����+ø��g��9={�ܞ���0��%�y����h(�X�ɣ���*��/���#�f ��������]�h��%�H	0ٸL�P�ޜ�_,ׯY��N���Yy�F�����p����Pa��?�W����K,���?��F4o��Ӂ���1�&�g�#E�*�@�9ū��z�Q$�HE�|�:�qhz���3 ���V����>�X2��;8�������R�h���G��	ɡnylOKoAz�����׸�ke���q�<z����o}S�CL%�Ρ�
�T�,�]K���<'�?��xѽ����O!�x�o=��쀬(Z��L����h��t��P�%�;E����2����^��ML�6�y�tcaN�`�4Q���_��u�؛�=���_	�av㇙�ڍ�q�/F��}���ג�6�wB;��ʼ�N���G�'.����;�[�J�&I�q�zu^���]PPV�LA!d�ѫ�V�\c_~;����L���=��F��VYi����kz�Md��Mҭ�3V���~gq+�f�o�O�"�\Z��,�%��|s�L�tff��w��"i��7��Ӥnp���Ǟ#����q��a^9���S�y^I~��13OAU�r�1��L~,���"</��	��ׯ�^��
���]�ZK<E�����x@��#܆�����:���R^����]KW[˴ew�J�Ǥ�y5�����J��0q���^���5ۿJ��q-_������S�3W?6�(��|b����e|����ܹ#�}Q㬅���aL^�r��Z���}lC�ձ���zֽ�\ْa�8
�T���~�q���N`ߕ��&y���UJ@Mj����X��)e/>#���L��P�{콅\��C�I�n:5�s���c�mZ�2vNb����#�$[	Vx��.Rt�]�0���z,��R��$T�p�y��e{B}����v��N%{Ӌv}�����)������Bfm�w�����N.�J��djdr9��"�~q�H�|�a�n����>���9 �+U��3%��0r:m��7����v%p���=�&�+)��*W�c�
�c=����}�֭�������@A���1�9�J�ӱE�Mm�)|�5�{:2y���oH=h��,����r���~@�N�w�uD�Vn�����OMQ�8�2r��6��nZ^�]Ly,��Dǯ<�C���j.3=�ݦC�}ҁڏ,�T@�k(�� �bA�%�0��n�|ayr;&g+{{����F��'v�������潿�^�NaRM��� �B�L��O�SLC���pA�����/����R %�����������-*�ωG7��e=���2�k%�~��D݊�~_i��a�o�T�3�m���э�۬�|O�lQ�f9��]x�F�
������NGW�O���o�R�|6^g'��opO3>�����a_Ue��{��n��;E�����8  ���]�JwwJI�=������^�b���=�<3{;4�~��Xjǧ�ߟ�ē��^�ը���5W�ʣ�4w�Ҹl��l1�0��[����zE�L2�$�vvO��At,+�㥯F�&u�C %xan4��V�[�%E���ibi�1���`&��ޅ�M|���z�����0����Ⲉ�O�s�z�]Ӈk4��� CmTQ�l�. !ۈLO"T�VE�0��2�s��G���vڴ�ܩ'@˅�����M՛Ag�x����б�B5�ь �ߊ�2L�<��?W#�t:G���<��s����;��<�����N|y��?ou�\"�7H�Q��*�1i	$�M��`�E�4M�/Ӣe"��>)Z,����D��%S��_>1���8�gS�xѽ�J;s���0o��ٱ�m�?��lS�5ߦ3P�pU/�ki2�465�{Mw6p�+x��/�+\��͔�tN�� G?����7!�w���PpO�ms����h����dPGT�h���	�*�+v��>����o	�|�VTz���BE�W|!��ߒs�¨���@_t�6��y=���3���G��,���ۉ1��>���+Fƈ�%e媷�tr<�yT�3jqx�h��˓JڴS�����
�4�������v<|��-��9G*��z��審���g׈x�;и���{�"�2�q�V"���e-.�B%�^F��Pf�*�f����
�o�Z�Q��L:Uwe��l������|�~E@¥�w�k�}K���X��xn�kWd_0U�2��
m��6v8���-�}!��R|��$����W9xU�����W�o��;'[rx:ó��sݕ��.בY�[�(������K������To�i�5��]lcP�qe$����i�ߌ,��f�X��
5��DC�¨�}�����gEU��r��5L,w]������M�l����3��| ��>Q��x�!Z�^�A4�Mdwa��Թ�ti�eJ���B�c��8���'ɽ���X䔻�U�r��s'��K*;3X���zkii�u;>���u'�5'���5;�9�H��.���/��{Q��,	���K7BKoy��m��q=��a��@>H>� _�W�츑�`�g�3%�뮞CΡK�B; ���1�t^t�=k��t���K��Q2���V.����HR6�(��(¥bʎ5���i���_��h�>*R�ף�؎������ț�MA�-�a��<Wـ��}i��m5�*�6�yk_w���+�zB����Q��q�m���=����v�q�Q�wG��p)@��7e$�����+?�5xV$Ю�=�Hg�v/'L9'������Sy$y�7��mZct��f4�����{�f��_�w'1I�,f��� eG���r ����ru�-E��.>/9�H>X>a~n��gL}���P��a�p�3$�2_b�(M<��8= VYF2��0�����ia����׺�B� [�r3��q�0Ψd���UQ��.�-�䫾�YX��^������"�	)�c�AP���di�M{�~g]7��W�Q�%Ʌr��pk�	���>����퀡�D��Ƨ�2*��-�"A����U��~�j����"Û$=���dM���ZU��^�1���ʣ��P���4�>���id��K�AGc8���[�w��B�#s�6��A'�Σ��I�%�ϗEpp����VՂ�M��An�v22��>�)����IMM}ފwq��&#������fC'�-��-���^���6��?��K�G�� V����q�7J$ݜ�΀{ ��'��K�ę�q；�+�|CnX�#N��;������EUk��.GM��}�X�V%�)zqw��Ìkm�C�u�+f㿥�=6�v����Fٯ۷�ñ��,9�30�9�[�g�`|�Ƿ�$<���d� �P4r:~�q`����Ҙt��f�����ӳI4H)�T��.�P6�O(��o ���2���H9��]IF����=�v�귍<�/�F��}kܨ�u��A�I��i�=�C��,(�H��M{ت-g�ˌ�py\ �I�n�t�|�6�-F�
���?[��?C�-��d��V>���WFG�mȥ��y�[�՞����п�!퇣�#Q����)��Ԕ"e;�����Q��?Npu�%�y@�ےP�v���0ޤ�g�탐��ʱ������v��px?�9vӵ��?���ۏ�҇ȇ���žS��{��3��xT�G�<�Bu~W��]��O��,�����ߌ.�A˔SMb*%����viq�Y5Ԕ�W����B�T�m���������[���yf�|���3`�͜%�7�/4#�g!�|T[��#��r��Qx�7�2�R����A��x��M�{�b�*�����%���>0�%~�O�-e���> b�P��qݷ=����|6��>.�rOzU!���g|���n;}U7=2��Y��z�X\��
�-7�g��'r�hfJו6�iP�M5���F�/�c�JOUw��� wXɡ&����J�`�˟���<��⫞Po�~;�1�N�N������q%A���(��b��]�W���Tmڬ�y��Rƅһ&y����i�
��6ѫF�ų��!5gÊ!��y��(�=�\�/?��T9o%ݏ��N�� [�$kr?s����i���L�ݾw�@���~��4yx��{5���ښh��3��x�[C=��VZ�zd���Cͺ�N���-���K~�l�Q\����4-U����4[���n7SN/�����w��&���|�4��`��*�]X�нcGN����%U5~bV��K�D�����Yr�ȏ��R�� Gj/�#�C���aD7����M�~���Ҋ5��R��ʜ�FQV�;k�v��΅0���Y�|11]i�z*Β�Z�� �l�v�tw&����R�Hɴ�kzJ,D�$T�[ג��3�Tԣ���HE�x	����PtJ̕W�&h~��:��E�]�,X���"�(�s��7�i�=?f�߄����IJ/� ~-���6Oh�}~aj���mʘ�#z�x _Y懦*ÈE�_$��%}�B<��vC���-�k�����0���\����1i����Q��>��z%�����i,��۰��*�7�>c]�d�}��g�ظǧN�2EDqA�)|g5K̜q\�^��	�P�ha.���O*���i^|�
e`�y�������Y&v�8yc=��E��1Б��r^e"�~u%���.+1v#���l?ʖ��z)�h�e��û����Q��l�kC�����l�5Ure!��(��{�6����	4���Y���V3ѳ���5{���D�Q���l״$ݟ��:�%J6����u��q�XU�1����Bt<�B�;jP*|t#Z�����D"��6���Y�w!d`n�h
S#1��j�:x\u�p�� wd�.7]��*��Ԓ"\�"�������;e���0��$�O�n��va��L�v�c�R�q27є��8����ݦ���������Gܴ���0��@�^2^4w��~�8��m��y4�δ�a ����b��$^����%
���f�1����r[�O�W���YHH��8��/i*�����IH��-�L�/��Z�]ɋι�-�Ԅ��0Z.;����RSI�ݏ��U܌vݜx�7�>�����m��� A�2
�U	�	5�V�G�^�T.�̂]�iHޓ������Rtk�I� \�9y~��9h���KwW�(=�4�
J�+fyL'�=[�j��[��]=�=�vh�(v�x�e�R�w���8�ߩ�ָ"�X%��5������N�&�yq��#�8 ��e���hKR۹��t3jlb�%�!�-8?�j��Uɋ���O�2a/_�KI��VG$.V�iTDE���7RTn�I���OsV����3�ϝ���g���jd�ξU�C�tرzK�H=�UÇ�jd�D�H�����Ib<_����\Z�n��)�i~��1{�Th���R@�#��� �8<4���a�=�~gt��-o<ȅB�
������K�=�k9�"�PV�R?}Q��ǋ���_���������~a�
��@2�} HS�{I���y����)��{T��O��5L��(_rr)2g��^<� ɑ����~�,ygN[D'$������9���'�Q���1����TX,�|�Lk�B�To�%��d}��_�&�dp�}䬼D*X��B��_F�v�zK��]R������Y��ae*ǎE���Q��i���=d�c� ��,*H�����M(�O�>���?!�L;�~�R-�_qߥ��`f�a���T�Z�� ���ȥ=�ܯud�K ��g_�-���?�&~��w����1D\[��Z�(@���O������)���'�p�WP��Dml�ѭ�l���>PPR���5��Ȃ;�x�+,Y>5���(l%�te�����4���?-$���zyݜ�W.��[��,���Q��]��j����[��$�́���f�Y�_�;�@�0p>w����yN 2��L��Xj�>��=�_
��ٍ���I��v-� ���W�|<�8�
�~df����n��h����a�JiQ�-Dh��5��O~ӫe"*�u� `f7D[�������(�Z=�5��{���

��M����s�������.-q�X�ggg<�S�vw�5hh]����3�u���K������ptś�놅��8��N��;^J(e*�������b'��z��y�y������jt��+QI��2/���I\�NSK�G$�>�RHJʾ7����/3S���'��[ƺ-���Q�Y�X��ar F�2�p�3�0�R�a�Q�(q�G	�/v�v�)~�Us�§d��k�c�zk9R��L��ށ�#GU}٩f�J����l� n�yHɒ�K�0祜\�	�%�W)�k�Y~�� _�uQ��q��f��_�������E)�Z��:����`^�$�����6�>�	��� v�>����6����r�������@GDN�tS���[UoF��N���b���-D�ڔA�PhXh���BC1_
CIe��E����p@��E�1"e���S�PI{�<�G?�a�(��x-p�0_F�AIE��d���>OC�B�f��r2��0Mql���/�C)� ^B�n�濮���x�`��r�L�e*7e�6�x��&��#��ňB���xi	����&$������q�7������,|��M�r��"9(� 2��mh�S��EX�rޕ����@�10�S������)h�����AQ�������WK���2۟]ȫ��H����$S*52�zb:��GL����S^�?��e�� ��O)0�]R�㥠�)>7L j���k�)��Xz�O_���@eP������M$w��4�S_��Ͳrc7�71�3\`�~á�gو���7���7YX%�ٽ�׋��] �"���u&T��ݚ���Y����ү�
���֜��Iu�i������U�M2�La͂�+�E����Z,�)�����Q3��������k���� ��a�<p����8bI 2f�bo���4�f����G*�����V�PN��".�ݥd�J�Z<���jV1���)LR�����>�"T�l�Ki�ϭ�T7��-G�>�XD�ԝ�ʆ/��̂͗��J�_[�w�6,n�9�_�y9��Ҩ����S�vF��!]�Ѫ5b(2ﰰ�SEU�SY3\����;e�Y+��v�����/�)	$���6>#��?8�/g#�b�]���W&-q��:p��M��ʩ?k�N�W"�z��gF��d)��?�`'�"�4rW"����痈������%����䌳��t�P��)�Y�҄9N��$%h	P�F����e�W~����6F�R�������'T9�;tC@0c�DFFh�鯙��Z�N���b��đn��[�i�q�V�D �;��?�Z4� I����Y��*+Y�TjIl>$c9�	���D-�}"��ڇ˒
?�����0�g��kQ�5l��S؀�W���
/��M�IYe���eo�qJt� lF"��T �
�c�&�#��d��4O��e������Q�5���k���d�9�&)/��a�Cw7����|��M���?�N���� ��%��Hd�-�����.p=�0�,�|��T�#��Zh�_���U5��E~N�ޟ�6�ޒ��,XDA���_�S�i)?VB��X+�.l4���Hv��^K>�+���Q>S��@=ߵ�&�&����k��:�
��.�VGH�з�'�r�qJ�$tJ���/��i'Y��]����]�p�[��_����,��/H9 ��exY�L윆���０���>*cz��n�~5��4 �쎭�~��i�f�4kǕ�;�(ˑ���m���/�7��u�ߙ�F#k��i�Q��Z��md�&X��
�Ѽz?-�2���Z�<a�� ����3���cc�|0.*؜(f����Qb���I7LOiT$����13�����mA����MQ�k6L�k��,��)���^�x�����5�:�rU����h^q�}*p�Q�mK��v�	6��1V?�����������>X_E��G"Mpb#�ˮOC��j�4�{�X�L�FѶ�Op���^�T�=)���I�-PX@���0�HU�.�k�v�(�~<3��W"VAo���Zk�%�Ȅ+��K�+�1G�x�Y(A/:t���c�(�~ΐ+�&p�ha�*��]R�k�+[}����[��v���������D����OШP�1�~��#	��I�ڴ�e�p�^7�p�C�;қm׏�!�v�h{<�A���(�����1��n+�b�"jց��@$����oE[N��YJme�Ax�>�	�a����|�$��f��J��'˛@�WV"�Nd2Z�*�deb�hH�xh�,f�G��B�����u	��O�K��dh�0��<嗗U�7Vz�	���n?łF�a�$����B7Dl�ds�	ʠw����z��Trn��
w��l��ݡ�������P,��&���c�!����,�;!f�"����W����;%|԰l�@oTd����7��D�����h�	f�,:U?g�XM���m���s��ƫl�/����:�.�U��`���cD1+�.��(��͠��o�#���� �S�B��p,R���$��Ri̹�)�>��]����5�M�I�>f�"�G�z��l~.�aJ��cz��3�R�|�߳U�3_N�$�&C���-� �4C�y����D:����v��]D�������2�l�4�\���[7������J��Z_W��~rG�\P�;;"՟Q1pt�ؘ�ѡ5�{������z?Y���"��uj]xUM��=%�6W9��?�� ){��y��A�P������ۊ���^��!t�[D"z�D&哂���OJOW���wc7`T�`��������FO��b�e��~zwED��d_&꠆���������w�(���õ-����=�����˷��h����wye�������J`��s�%�/�¬�"��vO÷M��Fy/��׋|x���$`��P�t�! ����XN
�U����+��{������؉�H��� ����^�긆���v�M�\]M���"d��9��we#�p�A��36TV�W��ː ��2d����<��D���T徟n�m����}D΅�Y彑.)gh|��vCs���pF��+��\���?W��9��T��e&�4%5��Z��f���
�Lf��#D
��"$�r�����=��O����|u��(��MS�Q�gW��㖚�߮�E���k�z�:k�c֯G?�o�?��K��鍟�2,�����='Gj|�A<@��~�|O�����P��?�޵�|J_�f�M�ڋ𯟍��Ip©�I��y�����f����}�>�e�\.|��u���mz� ,'�ۙ߷�AV� �[� 对��뙹c�J�m)ÙĔ.��9A�f�B���̮����^��d����[)ԁ�T��c���%N�MqI߇4����=�R�mUt��g���6���u�a�څ}�+jZC{5D͎�ꗪ��i��J7Ŋ���"�GYm��c¶��jn./x^�H���5��Ѫ�2���	§�h�����Z�m�cD�5� x�]����r���c�D�>�/�!�H���_��tr"��Ռ��������'���#׳S U
n���؇�ܠ�"�q^-�G(���nE.tnoP������v�	-?��������2��r������B(��{��'g�>W���:�V;G��F۲U�=�r��a��km&�	nӜ�)��ᑴ1�dZ�	U��
N�0p�Ѿ��.q~�$jM-�L<�Y���P!Q>������]s��4���v��?]΍_<5\�i���S��˅RÞ���g�сL�ˋ~���˲�	�]�Ǳ����	ײ.��ݸ�{"�݄��|��!�ْ��B��z�L��"d��,VBh�ևYC�;:^|�fv���^T��s帪����W@�������ɲ��t9�ǥM�V�΅݇(��\Ϋv�c��X����m�J�KjN�idG��3l�DE5��-��~e�'}gɒ��VY�qư�G"�e���e�㼗eKYV��Tv�{�a/ө��h���^�|�\;jC5iM�i�h���j�?=k�N����Vu^ko�� �d̙���w��		�q�(��<�ׂ����ߔek�*�M/Z��Ǹ�U����K�ʄ��7��y}��� ���N\':m�����ll���6��)���E��eaҧf�}#����Cb����ٝ2(<4u;��Y?O�Qf�r|�Q��nRF�X��jţDe�Vs���T��bg�ƚ9�'�S���ݔ�v���8KAT�a��ê�УC�^�!h�ytڙ�p�֠+�LXL>�Y��I<I��4g]���,�O��O-����F�js�`�X�9��0�mz�sD_d�a�M�N����&�����\O`;/�^,��P��J�FH��RT�P)<��0��лMg���Z����=_�U�|Eu�~
ٖs��f��&efu<h6�1�ɛ�0Ϊ�� ��"0��tfk>�\�Ys���^'�퓌Tю�z{���d�}��uͣ����h� A ��-l M�!�_��Jv����̒�
ϔu��6�ں/��k����RxMtlw7?R$��Iy�Ǔ#���]��
)�YH��b�R����֜��0"ݕjÍ�r��Q�a�`WR��?Ķ5q�yM��O[��E��M��r���,� �z�R�J`j���x��e7��ݯ��!�����}?ڻ0"���P�f��+1V��ξ�3�����y��|���qI���|�_z���e��g�4�(�F<�Cr����:�Fm?��:F_.'DvO�Z2*kί�}@�� ���� $9��Ȕ1��t�m?T���5v��gu'Np����H�ÚU�X
^n� T���`Ѧ�eLA��1N�X�օf����>�ٛ�dQ�iO�k�l_�1:�Rȶ�;i�^�p3þoT�_��C@�7�P����h�(�u'�^�3�r\*������$�O逽D�ڊ����'�F�"8j��,�@�I9 �OPM��	����ݠ{�oȓ� �?]Ǟ��܎�Gf؄S�Z�~͡����7>�d�k���h��Zm�W�j��V����@�)oIQD99�[ґxNB�� sI�~�����Am��,��+!���|��?)��>�0�_���	G��M�I�{+G̔�u#�����$KH��d\��]Z݂��rΙ����J��!V��ap�-_�<���]b��P�{�4:ϓ���]������M\��U|��rt�e ��	����� F��S)Za���ݱ�7΅�ֆ$��N��]+��M}�T�?J�\��7YA:�v8"�>�EE�z�=���|r^U�����7Ŵ%1��h6Nֻ��`�i�O����c�P���� ;�m\�P�m� �ٛ�G�;��ϚM��OLF�k��/���q)u���2z�9��B��_]W���M!K������k��B�c�3m��@�E$s��p��H�}��iZkSZ�F10��-Z��5y�J�������G&� ���I���� ����Λ�������=�Rӌ��M�C��n?)w<�p.lE�`���~�	�"|�`lԷg֡��,5u�^� a҂G�8�c-/Wؼ�B�G��"C���,���|,���z��V��T�oLS�qT��0����c@	f($��	v�0Ć����� *����2�&����~�1���2=��3`���H�r��Fv�yO��}-	�}%�{��%�M�d�KgD�.�Wb�b?4>��/��7��J��-����"�jR�Z��4�5_g$^ˎCo�{����+��5�t5�g�8�r��UĜ�
x0hI��Oߠ�:��@ff���B�E�������9���t���3�y��VB\f�w��ll�k^ӴooOW�J ���[,+8=���8V��CY�'�dW��;���z>~:�,�Ua�\���(�E^Y"��9�{�`:��?n��ǯ�)&�G���_�wE��'��Q��9m��=�ʇˢ,--T��>�����a�_��3l5@�U��Ö%pU�/l	�G��E�ϧ�=�LZ����lx��wRN<�&i��AN�XjoW��m�@������m�{���PՄ5���4a�`
d��xg����;?�FU\6�nTk�H%	���Ɣ��1/�:_����V�Sw��u�R�4�*�� �K^ �q��y���)=�/\1�	R�g�׃$w���!�$�X���Ӓ�eg�₁qqh�t2ye��GrC�=o��?�)�6���]jp�	к̅8�����
�T�/$m��u��y�g��ޓ��6��Il�nnp3lPP�k�f�d�	��s�rN���]��w�I�`6��/���&��l����[6�	������c���b��\bj�Q$�ڽ�|Ǡ2*�F*��k@j��VS�~�ss�^T1�6�|� R�.,��Oƣ�	�<M"�櫛����ΘC?��V1X����r��QA_���?9~�2n�[��]���}�b�zx�glp9���<i8>�.f�_ʠB1��fU"���&�	��4����JG�G��	E���
��b������y=iC�̱��C�3c��Cm�l�j���c�gL�a=�I��Xͷ�K��u#�ݗ�*Q�r=� �%C�����	�z�W�h��r�g�$��g��dvMbKW�^��ě(�T$Ό.�Ob߶,A�\o-���Q�2l�ϓ?�Y�;G�.�S�%������P���u��Z�r!�m�'D��B�ĺ�� �H�سy�سo�1mR��g�Kڋ��������qƏC-R�H���P�]q���^����qx`k��<�=H+b��Cf�0��h� �z0���$ 7��n�"9�*@�	�\����{
�ajv����Y�ns�����2��ae~ђ|����n
��+�`���.F%��I~$	��sń:�l�=�Up����[P���^U�cQ��� ;�[J���J����m�
���4  ��c��!���>����w��4�!i}��ihku�	��ƀ�B����,�ܨYpV�+b�."�Y�v���._ȗ��{���\s[Q����A���4eh5��O���[�{��m�~-�韢��s���vCh�4{���\y��v��p|kMSTE��1��^]��������HH
K ����5���.��F��n6s%Pv����b�t���i��ܪҾVCz��d�)��y��<E��7��,�c}���vc�����ᆎҎ9��x�}3��֌������}!	�$埏8ϧ�<���WS�4ZIiyxT�����rn�M�M�I��=Tε�����\*�����d���ԁ#v�d^�Sf��*�K�Ɂ�E�:�%��Q�Z/��~$�骒S~[�'�����������5&� .}~3oQL�K�+4�7s؆�XKE�Ν��?���E�a�E���2���E[%/�<g]���cm��-��"���ډ��I=k�V�\�%Z=�k�YɈ���W�$��_CQ�!���~3��/���.)ԿP��j� .�IG$��o�y:sl�*�<3YƦ�9?|��$��g�\�����G��:�o�6��/���$7@��w���ߪhfϳܸy��syLRY7��dwJ�_�x4�FӸ�至�t�{d�TY���?vC�e��ǰ��U��E	�N��P�i�+NQ\��t T�,�N]��5���L1ԯ� .�}E̜��n@���]���k�t���F\���3�?�RH��M������}<v�56�7�Y�jkC�h����
J�W���C8����"�<,���&�y��n,�ů`{�b-��{�ğ/�P~9���S����76xN���n���6�DP���D{z{ BG��`�h~�D �B�Q�x3 In�����3�\8mAAAE�)�ŷ��E��41��b.��/,~ᑄ5)��������Ld.|h������D��'A�����֑����c�9b#��k��r:��%D|Gg�qG3��7VF�C�e�͑������)�H������ק�n��zn�qI��gUsז�����ZHa�i��Ow��#�YH:��d�>����*.��kF%�`��y���Т� ����%v�J�Oǣ�*�����K��h)������T6Uzq�ۖ^��I[0� ���XaF��&�G}�8�!�s]u��h�^�md���w�Mr�T,!��@��Ǖ���t��]�x��gQŇRX���o0`^+F�Pk&��pk�Ɖ9%K$P������@�Γ��s7Q	�w��h�e��r����̾|���zb�0+[Y`r콻�E�[Ф�zC�]�3+y��=1��D�P��l��j�G k*����_Q��""
�_��i| �b���Dw��������� �-(�h��R�1wnZ^��"Z|$��EI��	r�N��y�QM)�H�~�(vr�쫻�a����kd ^�&^�~-�!�YZ`n� �P�T�w�A��@�Y.��m�č#��2`/�3�f��{�#Ǭn�����w��T�P	�	k���!B���)>@�.u}>c�� -�����)R�)f��o׳5괝&L�	�]>SB�z^���&Rvv������"Q�w=6F=}rs�$�����4��_Ҝ��<\f���1|J���MhI�{RH4�|�d�G9śj~�M̦vn]WCLH��0��k�b�Ih6��W鎂��J�Z���J�!@��gfd���ZpU��T���>R���i-.�-���U7_0�?MO-E4���8�$�6��Bެf�l?�:�9E��*{g�:B������鈞��d�Rޘ�@���=�V�(�N<��>k:�h+�C�w���!�؊�i
|�KEY{w�~���~���J�u}ðǑ���d�M��c��?T�)�l{(N{z�`�[�^�EE��{+\D+��=2���l?��S3�H*.1�S��Bq3���YuMS<c�@��osJ���sQk��$�W�.l�����E�@
y]_��)B�)v�� G�hm}��K%���l�yO��;h#��܆�#�$#�����<�ҫ����{?z���V�8�7�z�^��f�:|��2!�GT�r���D�*���](umT)���)�{��#n�H�d8c`Ƿ^A-�~�ڞ�� �R�7�gfI�lC6��Iʹ�{�ޓ));����"����+k������j�J�2i	8<$ �ƫ�f��)��k�˛�uu�+�~��uA�E{�_XP#ZPGh� 2{��~O�}����I�*��4�v��#�r����Ǒ��Q ϣ+��*i�$�#@��A��JV}��DRH�[�wMR�Y[1߷���>88�~_��ʲ�����\~�@[�������	J)w/��������ԶQ#��$�+�������U<#&yk�}��G���E%o@�t���T]��|?���Ra	��[ICD8{�"�������V���}�e�c3G�����I��e�hebL4:�;���?%7{4,���ěh(J햔č��s�=Hб����m����'��1���_n)+�ƕ�F�����h�Uи�����'�z{H�-}�!��"91ܗo�9����E �i����.%��a�1��.�q@�s] �p;VB Dkqq���
�c�1��ܼf煉��� �������C�����|��6mL�Z�&������Kީ���.����X�=�&��aǶRj����F�U%�XI��dE��J�EE��C3濓9-l�������PaO^R� 2%��l4TE'�b�WGik(�X������L4���xO�S�r)���?���v��?]��\���(Y��3}�}�:�9�sW���G~0�����Ǿ�R�n�x�8)>�0�{����%��NQ��c��^D���:a���D|���*6V)���U�#:�a k��.~�|�������=ooE��7�U.t�>Ka?�`yu����>�p�֥G�����|�[�6ϋ��B񉲾D�grZk���� �s�Y�����ٞSS��+�k�f�4�}���������P?3��Ke��^JbB$�!���R˹�IW�ڬ����x�0+�`�?_
�;&餝��:�0՘ɘ�38h�Hu�ϝ�K��7��h�
���7�֝H���rL֛@���3*������v8�>�AL6l����*��UgR��!0��2J�D�~�ˉH��D9X]��#�|(��\&3��/��E��'�D�7�)�juV'�O�C}"��q���	�&�d�ft*W
#-r�K��&q���ڸ���B?�cD���2�1B�Y��W�3��K!��p*O�M�m<V�%*G�ڴ8�U2X�5�6j)] 
"��|�A���gdzu�|�y�J@�uZ��0~�?	����7Y<���;��b].�����k������{����W���;�>E5��3�/W<�E��R!�ś17�Lt���_|�ZU��,�`m�7���7خw��]^����.�';Q0��+�V���S�O���0u��迖T����҉a���Zxԗb�2��jVm�-Z����=���?]!�3L�a(�U]�N���6磩��s]ʼY�� ѯ�thU��y*�,�'��Á[	��xZf�E#��4��Ze"���'�L1�Y�&&}��i�����,�s]���JXM�r�1\G7O�&)��x��&�@�
�f�	烃͕X)���
#ٸ�˳F�ǽ
�ڢ���	S4�R1���*�EUy��~�ɂ2Ԅ����Vq;�G����RoR�RRm�M6��.��8̧:�~�0�6B�@I�n����6�"�� �a^=޹!w0F��܄� �q_4AF�a_���!Y�F�:���f��1��q@��<d�f�_�����"�s��VA6L�c�$7�C���R�aE����eK=+��;뎁ԗBK��ۃ�چوh���k���j�i�!�5E{�ݮ��K�����]{ID11�8�>�.��!T�-c㉱ƌ�7��K}�Fa���"sA��*"c�	��s��Q�ބ����j�j'1E�%6�Fps���89�.�S�#��0���f`$#�0��|���lj���cb�:����&_{�e#ԙ ��Rui��U�&�>��媏��-Xpu7�7�Wcե��&:tE�'�bl�/brG��E�˞�-: cQQ6�%��=�9O���Zk�@d�
����b~T����~t4�o-[l�E�,	� .��	gk�[�U°o�@�����lq&�Lo��+u֘ߪ<㤢��������Z�A�8J�
J��8��<j,� 3R45<W[W7[ס����5�  �����ҩ
Uѯ}B�;�ΐѬޔѼI\<�m�S���3{\@Jf�E�^V��
E���-O�f�
JN�O���UU�gj�B71�2�-�����:n��p�<��o��'`tw2�#�xB�]�z���� y	𘡓��	&U���^}��8�Ҭ�9�I�����à��A.�O,�Za�x�DE�^�K_2F�3�W�IL@Wf����_�6M�� ��W�|�h���s�'fx{��(7����1g|�B]���s4Q��츺踤U�9��_�3$~8-����2�������3�L�&mFu����[R�W��!���ܶ�r�f���?f}��{���Vg��+L�gۡ��x����W��̙/��2A_
-Fx����U~¯:�$�Q��P��X��Pq�'&�fx�+�Aν��rW�Ɏ�ح��c�z�e�[*Y���^AZ��d�KJ�x�� 5�Y=I��+((�Xp)�A�l��g��v���}Ʒ�9�_�h}�,�Xp�ڒ}g�Jn�X���z]�V�Nn�k�H�` 2,f1�nHIї]vS��Ğ""uܞn�~}�hbHpp��N!y}�2�+��rס�P�7��t1uv�7zBxWo�㍻�2�'/2Ą�r�}ؿ����KG�W����9b��p�#�Q��>�gO��c���9E}�ձ@�K�����."  ��KHjA� �B<���������@�S]lZ���_~6��FR�c'm�s���a c:�����~����Yqab=��~tH�Ј�n�*2��*�$H䰑qQ�h�S%��F=���R�����T���tմŒ�y��W��?�B":"z･��{'j�:F'��=z'�h��F�э�;c���������,��{�>{?�����f�'�N)~�(�U?Jb!=f$=,��h�Tx��a~�I�~`��[���|�W1��Yu�]������q��p�̦OJ�
�<A^Z��K�"k�Zkw�X�r^݄�5����?�Z���M�~�yVϚS9����Ph}�O�>W~�_ʖ��ץ��|gJoF�[��y1�y/D�M��)�nT�L���E�iB酀�C=�~O�6X��4h�����Ot�6~Ց�yo��Y:f�E���+E������n��L#��6��;��2բ�����{�	E�D`4Sej�U	��o�hC���ObN��Ub(��JD��������B-ߕ(���K�i�8j����>.u���䇮H���=O��o�ɹ�)j��á������I���NA��a�_���Wt�d@=A���o+�(
�Y��y�9������_]]���C0���܂̬�}����Ʈh2�.��{XP�iy��l+z�!⒉�m��˫C����	��y�џ���Op`�>�"�IGG8��x�?�����-�N�r�����<���#�-��$GZ�c�6+�����W��yk�F|�j��iaO�e�4TJ�B�~�������$��HK����3����~')<U?���%P����<��0�49�@Q��?E���T����D[��Ջ��X�s���b��F��S���Uax��v���k�T"p�-/R�Q)L���=w��G�4j��J�K��6-:@e�D�׻���Iģ\�,VG���1�ao{���#�Qz����߻'�6��O��<܍p&���QDC�*�3����o���u�
-Y�68�,�P�fR?��&�
S�������8�,��:/��Hn�2#�m���8}_���/u12�賓df��wa�Z���ku��{܋�������ԃ��nN���ibKY@�Ȝv��{w`%XB���?����t�涷�Q7�
�vUw��bJ�=Q�/z�ۈd!Vg%�4�vF�^bUާ3���M�fs�4�]�����a]�!RD���,���d��iEՃ��BG�I�{߆ku�{r��NN]4GKX��j�#�d��>�F�4Ӳ8�F/ׄ�2
�=Ff�ūN�2��kb�&��
S��y��N<��ڴO�Xq?	8�N�w'*~����jr���F�&J��MbT8�	�(޶��a��)B��Q
�jU���չ[�[��}�Nr���e��O��Y4T��]7� �Va���<���0�21�)��|�L'��'��R��i�*Pz4=��l���]�ZD��A㋦�x�@4��#'���9��g�`��J�~XZq5�x �D�����iB;�&}�	�Yh9)JX���Fl�Q��P"�B�gx�U����Zۉ�c��Qj,�R\	?	��������X�.C����x[���l�����Yv=�4��Jy�����c>��oهV�#�i�Bf&�>�
�)�:�\`��5���F^�&Y9�c }j*�g�9Y��@؊�=�B��Aٛܲ�yx�L�(�A���l�[�ңf���+��K�:����S�V9�ϒd�� G9�&Ed�j��+��^�v_7=�:nܧ���������B��D
����i�)����VaD��#��~4�-��+8�A�HM�s1�_�H\��#�V�F������SIl�E�;�s����pu�~�ɕ�Y�~9��ӄ�4��X��C�f^�Q���e'���9:엱�����|"_ʉQ��<G�*�Q�'�"��N]�"F��}��'mD�� k�Y����}���(C4�3�����������������r��sM�-�\21H�,D�A��F)5��p�C������)/��迶>e	��>�hv|Sj�{�GA5��y�ݝ�bU򚟳�Hk#�{��̗h��|�<Q��_]�{u��Zi1�@;��m	4���+C_(���[0��8���H7d
��Esd�D�ٯ����_�~{kv������i�-XC$
vg����r[����,�X���J>��X>=2�M�K&J���K*+��/���&��TyI���m��U��օrf��\j��m��'�,�|V!��b}�8h#�qY����9����fb��@��w�yy�o!b����S�%��s�#��V�!AKY#s�'�Z]� Ϸ��K��T1��gE��nZd!h�JA �E�p��:�����^��k*U���ia6�%Y��3�s��R�-����v� ���������{U'#_V��.2��Z�Ļ��wbrJ2��.�����j�ה��H������ą�����c^���U�ݲVpP��S�	�0��/=���|��K��%���/Ŧ�+Ob�ښ��	�Gx4.>#�����N��QQ�y���yhհ��F_�i~$|(��_�F.ǈ��J�%��5cAj+��8�t5�N46���A� UXگO,�@�}oSQ��.�������9��̈́�Y@�b�ݮ"t;���4r��/li�*6V���=����v,�|�9���f��Vnr�+h3��&���|k�Qi�E��F�%1���YRV6B�,��¸�w�N��S��Z�kV�$��b��ⶋ�\jMp_��=���S��0���m��v�GЗ�~̪&?������g_��/ui2�{��TpM�k����'W��9K���V��/޴�Z!�	fjĤPҔ�I�M�^�AyG��!�{h���lg���ǻx��=����Z����hE�X�	{���K��3��+ėc�����y<Q�80������)O /..>>#PVs���\�c�ss>͘�����A�,n\�V{o$��ս��6-�{��|
+}�zq�!�tG�w$��0��甛vטK�����n|�����e���ٲ\�ذr��֝du�]�a�>�ه_ˡ%mרf��-���g51vcK.(��:n4�Ķ�T} ]�<�L?�S��G�Y�>C��W�o&�\6�h����ū��|���n�x�_���-�~Y��{jz#a���M85V�M
A�vƦa�7�GV���w�+#7��BϨ%/)�F#�U�৘�qjO�߾����u��5B�g)/�ߞ[�X���[��xtUᐔ[�����Ϸ2��י� �V�u�-@[���nC����[����sӪ2�ohf��Don��59�N�������	�[:���#Wv�a���5����J��V�5Mڰ�2��0ۮ�k#�ߐ�w��J�\��s= ����n������(Q�$��b�/v����P��ς��DD	^�����\9G���/���������g��!� N� sao�����#�7��u}��2�#7:]O�SWۡ�홓�m�ߩ����|�J�H^�1r��x֍�'��h�?v��LX�f�*�:�˛7K���Ø> j7��v�jY�s���M>���Ksbt��[۪KQV��.��7�'~�h"	�������̈́��hG�%��4[>W�"��K�ب�h]RS�O�P�;�Λ�<A��I>�yo}H�E~��fC�JC�F!-��_��f/�	P*1)n��!���8��� ����5�ԣtp���B�<����J�qui�k}��m,䭋.�<ڢ��@��Խ�L^n��&��;�9w�-om�ޮd��qj����)��W3�)r�+�SdK7iK����\ׅN�;�7|�D'YȬq�\��� 4C����-���1�n@����H��2�%��3�^u��:#kv�:�- m������-�ܐSV]��I�!�w�ш����g߸s9W!��d	�R��E̋�Z=�2f��}�������'!�;��\g��v�.����p�	�>r�#As4j�Lb��s9gr2}�?�8��8�7�I�}^������JyH` �_H<�Wqq^�ո;��x�a,������2�L��m���rAk�
���j^��r3��`#Y%2Y),o��"�����
2�>����_�A�����Qui*P|�4v�d�t�/:&���T�f��G�<"V�=\Z9�d���A�.~t�z�z�3�&8$�4(��|�,��FT�fĴp���D_�.6L5C[�gOҊ�[|��mIY�`�ݔ9~�}«+q�6�24���O��cpH)��]¤��R[�B}�~n�n��C�����9~���V�Q���]#�b���S�;c�R�3X��nk��ѧ.+t�4EHg}���^�{���׋�p�*�d���ݼ���xQ��.��Ï�:#�2��I�����z����Y�q���I%�c�zt���1B{�6ވ۹$Ew�/���6#�j��e�j�t�j��Q��Sd��ɗ�V�$�q#��E�Y�?[����W�ɲ����}H��Yܶ�頥�ؾMc(�Զ��Xk�2?}X叕�z�q _]r�%�0�.�lƶ@C���.Tz��]fV�-k�Gr>'$�PSfDg�:�=O��2H���WA�#=�>F�dv��.� )���w���{�;�6��\����s5Α�p��ptd-r���vcֹ]�f���?~?�;{����4�\7�5U8i%L�\�_�ڰ���jHI�vY!���6��أoО�����uu@J�ծ�z ��V��1���wZ��@0l�B�����da�����% /���-���l=���=~�Уw�^
a0��\��O�o��iC����.���gj���[o������J��m���
%s�留�J�n�� -�����{�֟
.�Q� �b0��ڧǈ"�|���錠�����٭1�t�CاT�C�%�2�ވ�oq8 M��e�3sJ����O䢺�~7=wwc���� ��9�ݴꄌ���B=_�?���L.ڨ%�/f	s�"ZY�'��I��c�������	O���r�o��nd���xF�fJ-*�������vMW�8�q
�~C-諪]k�4�����+�+g��'������<��^��?Si!�J��sz)�]�=�iى��(��6 z�{d�@��u�'WO�q�R��_|�X����n/�I)�p�
��A�]����"P  ��U_��60e�,"�g��������H��]~��:�hS�$�nm?��� ^�ؗNy��6`���芶.���;���2ܩڒ��wC�2�t.��1f	��l{�Yه�G�bsS���ێ���٣D�o�~���p8��!�~�b�Q�wG��nn��du%U��+�4��4�*	օ�f*a�9��j#�!��ܽz�`L�l':-a�k�NC��Z�:�.)m��5/�����4��%،��k+��[�޾�G�Ӌ4��wѹϑ}V\�����߈�o1U/��1�Zo����>�AW���(�/3$7$J�&a,=���F�6��J�*�bB/�����H�<a�]��t�^-W�n�4��7����lwFDͤ��xZ ׍ ��@U�˄��z�(C'�J��Q)E҄,����ǐ�/�.����M���w��{���w���y��D̓F2�C��ܺ�p9�%h�=��֋������Ulu��D%��mh�v�)u�i�XT*3>N����D����_�\W�= �]?x���š��~x:�[�{w����=1ߞJ����Vբ��<�-�\u�q^�k��¥M	#�����'E��Ы��g�j�fI	g�3��Ԫ$Z�w�����Y?�*)�o���/�>��e������PJ�(
���o_q�����(����90PgiJ��h��W��j	��I��\���	>L��D������*լO������ݯ�y��U���*���k�R���h�e��GR�m7k8$6�H#J�S���!�z���5ėQ;����"����U���zX�o�ױ�),���U�ɑcf֬�N=u?6�(�� �zm�����2_��LH+W__��Ý��2�W��wE��H i�C}�s8;h>����v�|%�(���V8[���w��	��& �w. ����?r�͵� pT����Y���2���͏LP��3�F�q�k��H��^��Ûf���q}C}���%QH_Fg��,��s�Ӝ	�G;���w��������_W�Y<��6�e���(�=�<nӳ1XϬtaQiY�iC����8Iۻ��~�vo��w���ꍵq�{t���Ĩ��A������N��9���\�#���cp:���f���~%�>�����.���e��Q�䲗�E5��A[k<V�f/(��a���9mp��y�"�eS�?e���_�n�2�X�=�.�C��ka�r`�Cfw޺��X��թ(�Rߛ�/62%�"ӀO��
��}�=� 5pA�v�0S�6R������=�k��p��Z�P�{��(�Xz�b���w��-4��ru�P��r�j����\ٝ��E���>Ϭy���dJ-יm�~z�M�H��g�/5���_pA�kVN}^�2����'��/����
�W��#�x�H�-mq1S�[�exl�����[�����^m��v��%���ީ2r�@x�/<�bw��&�8��F�׈ƀ""�*�pi�C)�W��w�=D�}m��0�l���[E���r,�Q�4�.+o�1���L8�A�c?ǲ�dg�&�QA��g�*��ReD �~tuW$F:�;�4�f��s61�k
�������N�T��S�S�����Z��*f��G����L��Z˒�v��[`�\��J��|%����ͼ暰����7����Y2$�/?�1o0c��y̒g.��R~�D��@7�P2�:��U����T�w�,֪[���cbQ�w�/(Pf\�ú��RJ@�E��㈈m��BfjVX�Ԙ��?�L{�:<��x���u��%c�lT�!�<a�x��;v�o0����1+�5PBv�6��k����sB�����WS�"N��f#'�/��Dq��5��O �}��d����4�K�x�DՌ����G�\��ɺ߸h.{�h�;N�ǵ�{�Y�w����;���kB�:�~a|�@�ي��Kۥ�b��pF������BqO��5P{�����<fC�����xf<����؞���HteCݛVo�0����x��"��|e��hT�]P(�/���,�X�;9�
���`��!��F��ړ�dIf{Ǣ���Ӵȿ7�h��"Z�����f��u3�)9H	!I��D�R'�����a�d���Ѿ�"aar�bsk��8�[��\�Mq3Ax�=�(��� eq*�qq��R��d6st�q���son5'��5�oRZ����a1�n�����i,�zA#ã-Pձ[M���"�.AL�m2D��~�	�R�k�	;o<Z%��[sK�d��?|��Qx�Q�\���.X����b�;�u����
��z���/���M�uۦ{ө��Z�3�nos�(��x�,��$����^..q��:�x� �OFW�xS��.�ަ��{���tP��`�l���{��ĘY����M/צ.�^&���qG��W�1����WdL��ぺޒT�c$�:�׏	�"�NX������	 -��~�����k�g^?�Rx-�C��C$5�!����RV+�-�2����7/ �3���݄�1%h�ؐ{8>����{w�Q`�-�}��һ'E�&r�h�ʳ��B/�3�.��#����ȧ�Z!30����@�:��"&����mo[ʸJ{O�(���_��V��T���{~-���%oc�g�9ea��II�.ovm��X?R�~�3����	>���"�~��Gʣp�Q�}����c�@�����˅V<�ڷNz�V� ��h{R5#��2����&ǆ�P�ү�^I�����d6�� Xx����TFm���D���1�}��qF��(�A@��Ge6�n�8��x��@�u	E�~'���}�ܮ���U��,���v3��}�	
����g#�����8J�(��j�e�6�ɶ��Դ;�G�aվ�m5]P�O��H����;���R��O7s�Z4��������ٱU���|�6[
{�&��n�-�βP��```+%������+u'���8��@�(�4k���?���-�J����w�d<ZyW���\2��@�3��/F�ڍd�&�3��XO��s}-i��X����ϭm߆�O��D��O����?��1�Nk*���.e�-����k˿;2>�`�H�Km������������k��ɀ�������r��������m��ߟۆ����Q�	d�jkXgԇǼ悼�J~!�w��ˣ���?��6��]�'�xuݍ�=,*�6̒���D2����UX�W����<(矕�ϼ�o�ꇩ)c�K�4P����Ѩm��M�W���m"c�&)���m|M>�:��f���Un�/1y�j�(5����-�y#YkV1<:�ΰ3֙j�����Z��R��NL� �C7M���g�N��p2eC�d���~��gQr@d�fdť��r���ǰ�����$WnZ7���[m$G�����\����.s���{�@j�*B��H�\���"��2֥�*���І��/�#�rl(�_���"PU�k5�u��$_@����P��aMa[�%Q�=uw�>�ąR����o<���'��D!ꉋ/����s��I9�S�e̬K@���y {�Q>:�I�����Ll�:��1ȭ̆t�=e�_o�--͞��Hd�s�3Ӎ�h��"a��G���8�*��om����t���G����k7��M(���+ss�3"A����7��d�0� �q���/;#��D����	��d@V"ѫ[�O��r��-`u�A�,���W�,�����'��������s���f��Ҹ�}U��g�5Օ�R�-��3do��P����*��q��;�kӸbGr7�Dv	��㏃�F�-1�w;�!x�� H�]����(;MCy�L	P�N��y�|�8>�	�\F�=�r3���~� l��
�f�i������"U��^��@}�+���0h�YG?X|��T��"��w.bW�����q��:TQ_yC��Wp�\Ȁ��΀��m& ���މ�r��飶1�Y�I�T� :���\U�ٺ>�Bn�W����/�#��qc����=�E�=CD�=ϼ��J���+�]V�!�gs�_�T����Fֹ3�MPA�R�g�U�֕��Gm�����4V[5�zS�,��V��QF�PFM�s�_��3�F9�r���\~%��+����w��)*����Ok���j֏�>5q�*2V��K�>�r@��j��"��W#�cɆVyzc�"�~�3OW��i�H��M)T�P(גuѥDp/s�Ɛ�[g��TO6�{���$�Uk#v)��Q����])��4�"��٬���8�Z�S����e����V�F�	�B�=Q�p����v��x�h����|v��t������U?SZL�����2x��X��>�.X���J��7�Q�M��P��V���ce���?-3k������SI�~�q�@C9]������0в�Ț�IB"�w�������.i���i-�V�.r�ٜa���"|��8>�(gӎ��3��*O5J(�5�27�<Q���@+�yK��k6
�l1E�X���s�esݖ�/w�e��w�W[�v7	� ��:��!���q�e��+�
��s�~�ߞ'��.�u
t!���G"�	ZL3Ac��L4�z-��6��n&H�^�,Lj]�:��g#�x�O�i+�*��~.�I!g�v�O��P}�����~�͸��>�x���W�"��eߩUI���+\��K�_�����^�����w%�^4Iji��>T�U͒x/M�i�|�����!��2퇿[��!�}E�~�Zg�e��
��	b[����+��F��-��m���A����I�O/r�b9/�{\��Lt��#���G��Ϸ�n������M�n�1�P��i�m���'��aP˄���abb��ml�>`v��)Q�j2LO�q��t�#d�`��-��iBh����?�j"�rB��ŀ� �m<��<v���}fV5���DlI��!��V��:�-0{��iM�$��/���q7��TI�Ox�j�#�����;b7�KA��̾�w��c��o��y(�U���l�ڜ���ߛi���B�<ݦH�eY�����z���[Q��D�6�H��7Y�Ț�k��*��΍�E�8�}O������Ӵz�����뛂�������'A��0���UZ�+w���`�\ l�B;�_7Su������ R�'��Yd���#���ҟ7��d�ˎ���S�\�m �}/�ܽ���OC���L�2%�.��\�[��\��u���֎3Q�a�{i�+�u(��WΙ�E��n��m�3��o���i�ѥq��	�i�@Ni�3�D;��t�y�T�Dx�r��X�z��궿XI�.��X���o�Ea��[���'@�)<O�m�'4�uuQT�H�h_�0�NL8(�6�oFEO�^���v��LrWz�@w�.L�]tQ�߳��J^˙|����߭�}���F�x�#>C��/P�2��b�fq:��������m��W݈c��4�M;uy��g��fڵ�L�����qUc�+ʨ�u�[���5�^�{��2'{=��F���-w��ȟ�[S���?_��{!$�YO�	���
i^��'wu�x�&���0�{���D�&�Uϱ0d3s	�sh�LV���G�ˉ��8�A�j�#�gu0P�T���'���U��T��ԞY�l'�.4���������� Iv�=���S'v7.���&���z�ٽu-�:.z�+��\����n���D�''B@�{ŧp2�9ם7���Q8�E�µ�DQ|�bxu�����a�L~Q{�RM�1�@J;�nw��xgcGDu"���)���ٷ��c�7���ҙ�`�sQu�2X��um�S��@�	M9��K��뚭)l͓��P䯙{`j�����9�c��G=��^�9��Ʈ��~���Ɇ��y}QTeM����d�t�VdI	����R�dX�j9�V�_��b����WǵE�Z���s��׼׳Nt0�L�2fnu\@Vր����W/�r�ӻ��_)}���\/˻1+ۙ8;I�Գ�v:ek٨�ZK�'���rN��,����DȒ�꥛��}	x�����*O��V�k ��s�>����M9�'���ć����ԁ%5�HT�S�cB�$E����N�|��ü�.k���n�;]��	ӋwY��Qv�7R���tB���k;�N6^--��w�<��~)�n�+��(K8f�_+C���T�����Yن1v����c�儂�m��$mBx���ՃΧM�I��שٴ3DT1��Lx+c�� {�߲oZ�W[U

�gʨ3̄�r��������mS�,��#��t�zd*�s`���S�Y����~Z�|�x���t�Λqj��%���Y^Ԛ��2�,h��o��#��8ϸl��x��	 G^�T�e9Q����0�L]+� ��1���g�H��"���N=|���o�"c5�bWڞs���G�e,�O�)�.��J�J���N��mA����6���J�9������Qr��Mߩ|<�3�O�fw�C����`�g��ӭ&���Q6νv^_:a.Z�\�۞�{��.w�{b'՟XT=�^��Ak�Ϫ�����w[��s\F�"���^���󺀒��=ҳps�Zs�Ȧ��p�=�xE���B%��\pSY��5\7T�@�+N�de��a�D_�3��鹁�����ujb����7�fvE��!�����M����j����b01��i�)^�F�Lk�w�C�0%��2P�\Ժ���tv̦�PfYF���0u	b?�$
��2�yJFN�N@{���Č��#m��+{bÔ�H ���ym,e�|�\��Zp�H@�\�!�ztޟ<���3����kͬ�����9E�	�i��ά�,�z-�����}���E38����9<v�eG/�Q�B�b	#�P+���aoD�뙳�iK*B��a�q���$W�*�g�_��j�W��{���"a�=�=����r�6��	��Yᚋ��a�,��+*�:�s4�ST����J��u���E"ΆNoj�И��k��%�����z��%����d����UA�g��m��糉P�2��<Z�)x��C!na�WW������3�D���b��q�v��;�nL�ە�F?��|[�4W��ĵ��Ը��5=7�i�ɠ;we��[	�l�2�?��AJ��9�G[Q�����+Dl|,�Dq��� :�5e-:�X��pmwgӭS�W�I��&�2|
J��KG���u9I���%���RV��1P��k��r8���Ϝ��Y��I-��L�C��Ǡ�����f&��a�U�+����R�&!ƻ��I~��JB槛��W��^�o}�sn� �t�2�?����7>�_���J���h;j�q�1����N��s�`?�Y{U�����o��\����(Ε��)�R3��֥ؒ��r*O���=U|�[D[ٶ(�޸�D�ִ��>�ԐDR�#�ǣbwoS'�s�^^�|'�,K/�Ӄ���np�KM��>���)����ToZ���� �Z� �zcO?�Y��Ni�r���[kY��rѼh,�'�b��P�F�[��L0R�����A��k����O{�;;8SS3�U͕�>>_�������OSL��y{F?ɪ-� 4i��3dLG"o�QP0P?\�=��3��md-p�Z�MD��f:A�����K����1*vu��N�C�mG4vr\|�f��n�Pw@4�����r[n����ݶF�wc16�<���p}X��f�07����  �)z�s�g*w�&쇚�κzK̺��
�O�C�|����*��I��-ݒ�fx�L�H�p�|�R�s�.[���V���d��E�gd��Ř�d�ͧAx��T-�{9h�O��7�ɩ��dO"��Z���Y�*k��c\�g|��u[	l�~�?-�/B��-��8)�sTw$W�ys�:ʊ�x-��q�����d}��٣n�GbN�iyw�t���cC�`��$�.�w����L�j�1���7O+[ڃW3��w�Bu�B�&��U7G�k�%��XC�
�Sx�l��	�z�ט��V����\�(��3����P�f�[A��k�1?�D�e�Wz}���
�2gf5M�G˘�/�'}�?0.��x����%/�e��㯠�9��ܚ��HhQ~�������ge�����8�A����O;~����H\�'��g^Pyl��7}5q�r�����:u��̲D�U��o��e���ƥ��Tw��KB��w�Q%O��Q��(��BA6Z5�����X( ���㫆�~?��4'�o�%Ҝ�|�ϗJ����#]�B�*�	�s�����fnI�*Q}��^�o:��
f�0v�E��w��?��3�	ڗ�'c	Fr}?}-��ɗ�h�.��܇(���R�mw!���+:��,���ӽ˩ѓ�u��h�P
��ܫ`��K�d���)~�З��=�P�Z�VͲ��s=��w�%�_���y��<�Q| yW(򾄮��T	_ra��L�e�7����z�[W#	l�־Zvq�\���{�x⧥XK�=���;�-�"�͖(~�?i�iո/���/W�{m��;Lm�f���d�H���Qh�o�4qG���ѽ�u��[�!Mm������l��:F����B�h�N�&�,�]�3lrq�"�kӹtl���K͹ܬ�9;)�@�V�졛<���h�I�}wB��gЅ�a�v�'c�%j�*��F�Ե��C�1|l����_��-���e���V�-����L��ѹ+�G�x�	>~�^�k9�ώ�����as��	�r��5?�Kpaٱ�����{+� _4`�t��~(u���B�&`�T��D�,�1^���ۏ�2я%nk�ᕕl@����WlFg���5�s.j8�b��<^T�a~�#���;�igO+�.x�i�u���"������c�+:z��G_ݰ�`�����K�Ai,��bZ=ik��)�_���5��la\||���&|C{�E�P����EU
ދqŎ�r`�%}�%�M`��+<��b�lI�׍
2)�[:Xv�i(�����L�v,���W����<���=#�Nt��:�o`d��L�?t⭸m�����:9�xs�F���Z��/�f��A��K����'�n&bUF���y"Pq����Y2����<y�{�ͭ�ziYڶe坟��-�[r��R��^S�m'�F�z�(*�{��������(du�ڴw���L+2�9�'#�Q�֙��k���S{�c�}�V�r�����c�pm���͉8�ƚ2����"���m��w>����U�j��U�-k��av�)�B�w>ݿ�}�>�Uux��Z-�r������2��O�� 0�K���)v#�i:��_\�C�;T~�A������;��,�����w`1dS�y����`���8\��3�,r��d���gP,�������8t_l�&����:`+7_!s���H8+�s�ej/"��!���r߆�ٷܶ�%$�����Cc4"e�kP�GW}q���񠦩�#~n��
<��;Ut��FLB�Hκ�Q�SW�}r��U��K�w��Ke	h���p�͎�ۧ59�n�\�r��A��"Uñ_n!��[����p�	�� A껞�ҏr�ǫ���3h_�}�Hg���o�޼��tC�3�
������;�.*���%��J����D^]n��j��N'�42I�+���>]X�AaSs�������)=OR��O�iR�?I��q���-�NS��|�>~�E��R�?�h���>���ۉ�|fd�F2!������s1��x�T���1ېA�z*%��>�>w�v/ ���<�O����.�m���A$�_��7�@M1�p���������vj�x��r�N���?:~y3ݙ��_��A%��e'���-�-���]���fC�}t��n�խ�g��v�ݢ�p��hdpv�@�T��'ꯎl+FzK?{��}��勅���v��o0j^�������,�&�>���HҐ�+B_-�x�dx��8ЃE�#�,���K
D�$�=���1���l�%��Q���K����8_��o�l�T$R`W��V�Ť'K�������W�O�"��kS��W��P��|���Łs/�e�݄T�f�j)pe�������׭>��������#�uo��m��qӭ빙Vݓ~t��3O5">��n6�i��"�qפx��ڨ�S��=!��=�ԝ��a����,��h���b�t�,Ry��� �o���O����T�:�u�Z$��6�~Ѡxgl���������$�=���{�7���OlV?{����������%��ٔC{���f*�b��
�B���3�����Y�HVȵ�dn�Z*�YYG��{Z��'�c�_j}��{:=Q/��{�i�ӳ/�6�a8U���?�QT��qQ�%��7?Z�̇��*�$��V�om(�Aip�J-�ݿt2W�B�J�� �I�g���q��Yx��y/�g���
F������
W�hb���.H��.�y�`����i��z4���&"bso�U�3bxg�O��4�W�ۚ�a��c���T����8nYbY�K}X����1M��s4�|&n�c`�sI`H����-�on��{��R0*�k���
�@�x�-#VX�ڟ�i����{�%��%�@:0�m�k��2aS|��,B�>C��~��~��
�C�	u.�������;H0��_z���j��Gk:�����4�f��1!���>+�G����Ҫ������$f���q��q���ur��{�./>��=��.X���V�ss@i�<3�qE	��H�(#-q!�W	�ğH��_YZ�d�p�|�q=^E��Q�S�]
�|"��F}/ZD�������h(��;&�R�&��ǘ���L�D�TgO��#=V!1�E6S������^������k�,h����߄�o>){�8S=zq��R�}=�Oxxz��3�Ln>��{a����넹��n��`q�ff1�M�'ր�1��-� ��o��Q�- ���VM��?��h����s~��r��h��(��%U�0T$a�����My	�&�!��?v�aȻ4 i��Ғ��B�?���f��b�������n��IӮ������AU�\^��[������aO���$�5�&~F�όi���F���5�[��Da�G����,��:�Q�{?��XsIj�U��_~��<�c�b�A�D�z�d�?���D&�Ū�^n0\͏fz���1<Y,/3O)�¦����˷aϐ����z�©xDX�#F���ctEX$,YRmRg���-��:�ѕcu�u��C�=V":�|�:�!�{z�Y��_�+c���"ҢI�=m�u��4?Y�n�sz��+�fF��b�g��
kmtT��^ Ouʄ���)%����f8�l{o���"�b�_����ل3��F�rվX5��[d88�����^�q��\%8�.���;`���%���p�>&��^ ��O��>��`��H�Di�+�J	$��4MgBy+J`vm�풻ho�����T{���l �n����6�U�<e"�������������-���λ_W�;�Q�H`|l\��f�S��βp�W�`���Ϋ�5}�"��K��8��`�XK5^�J�y�Ig��y��մ��x�Uo.�����)�PlVc��4���)�k���͞��lD�hX��X\��^zg��HRR���G�.�wm��*�dn>��()uҠ�Z�?�p^Rj��[���5u�aQu_w@���DB��Q@JJ�T�qh��$�����n������o����;�Z��a�G���B�'����h��2n�א%vk�D���v��1�� ���lΠ��d���d>޽�;��ڌTQ�2�<UEa~��ZҸ��{�{jg@��9����!�.HdK���a���A�U崷`1
=�~�=@!������D�>�����I��H�<���L}�T;��4����*@b�De�f7��f����̐��;x��<�
�lu�
�l3f#}�S�u�)�rYڽ́䕦qEz=�����TA&�"6^�Hbq�lɦ
E�Gj�)P�l�e����l�i�CP����Y�A֨\f���,��O���`RlX���%��!�=��t�~�1����x0� �/_^��`���o��-��]>��[ކ��H�T͛4�C�ӜB��+%]�	V�7+�(a�:e��nV�~PctF��HH��]
�Ꮀ�6�kx/��t����2�
?�	��ɩBp�j`��2)�5]8��p�����D�aK�e�"_���\hui�z���]]�҇U�Ӷ`!��c��N��f� !!����@{������(;��qs���Hc�S�8�g#��U4iY$��x��3�Px����GBzF���̳iS�xV���Fk�r�j��2B[]�����b�,I	�T
x.�Nh��~�tJz�lz�6�u4�D��^C�,��-D�����E��o�9'��Nv��ro�$ߊ]ZxL��`���9��jNW����ZC|8Y���3�wr'��2#�6(C֢�L�G�eŰ� �]�e�	nW�C������,.�'8rPy����B�`�
�("��k����r?y��q�â�Na���ހZ�{���x�G\��Dk�aM�I._��7�@�C���r�(����M�jp��(@��&��?7���Mp� 6�D&���`&e�65��IHT����jMo��X]C��x6��S۫�L�
�?Rݛ��0���f���u�?�ɫ�ժ�S�X�,�S���;}epp*:W�}�0l�E����dXM�̝� �x���KG���U^nX�pxO��:z�l�|�1�4}J>�+Y�P$x���(�@���줂�yy�1}Jᇱ�Cx8�NO�8Ѹnc��;a��7
���B�U�W��OX��JV$�t�)��E�3f��E���������/պ��}�/e$&�8p���b?���ׁN$����f<	��y� ���|^T��+�����w�l$���#�Y&�@�Y�Ц��S�w�RRh^R@\�z(ʓ��p��8ʢ�,ۮ�P�{F��>�H`� ��H�6��<,@"�?�盋.�/?:��@��ȷ�猒��� r��/o�П�JT��ۍD2��S��,�HX��UY���䒅�7ܬV�LL��M|B^j@1)U�����S`T��a�2�D�hh�Z@iQ���l���""���4dRl��h�X��SH1Y�X�řn�����?^���u�����S���L����?R �X,�7���Ǆ1�L���mS���\`=똰�0*}6t1�����Ήu��?��e�㨫J]�5�`ﷆD'T�/�U�Կ?��m��[l�1���' �T���1]gt�~���i?0�LF��&�o�v��ӝ��y>W�5��j����>��µ�
P�P��a���?Kh2�_�V�
n˦��C	� K}'0�(ؑ���v�@��&-�F��fpޤ�m���0N�Lf��+�w1tU�/��=q(A>��D�}���:`i�>5�P�|�!T
�-�Ћ	����yKo�7xT�����g�ܭi��Y�Ѣ!P�|���raj��``a�LW�����<��Ճ�/x���
~
������|+���L~���
��y//���$������Pn~5��&���NH��I�����_욿E+��:��O��Bi��'������L�'r����l��J�xZ��
��X��P<��A�+)���tV�(	���
�?��&8N�T-bEU�qc����B��i��g:�(�U熭�;�:�b�èk�#��k�L �v{x�< ؚٰG4i��:jj�Q�O������7%��_�d�kĹ°h~+���(�3��û�������/y>Ϡ�w�+��-8H�F����B��t��ޕi�_���pq�n�i��w�sm(������?R~=g�T�ل`���"h�$�B�6�۠"�J:��Z�CݧU�"uuˊk�<�/&�	-��l�%O����Ҫ6�|���'��ކ��*����jЌ2kc
�OF�N�4�#mEm��ܰ�N���U����լ�p���p�a�����Ku�����w%c��rH���~��_�e�P��r;y-��	�+͜�9�u˪ ��`����h쟋5f��	�g8�����o̤��n�h����I��N��U:��(vt�u\��W������������%���Y(�jD��b"P&� "U,C��k�W��RS��}E�a\EM��׵Έ��i�������Ms=8���π�����Kje��E��ǉ�".�$�l��	F<�F��V��k�V��o��Z��u�H��J�̞e��㥥���M���| �� E�p�D���;Ɋ)��ez^���ქ��G�~pOV9���M���Ie� R��1�S0M�������!I�o줼tVǪy�\�Z}S�|���v"C%��1Ns+�]B�X�I�;y���&5�pp������6��6��1���6u�8�t�6�c*P�I��>�˰zG�*���='�N�H1r�Q��|�C��,�G^�+�3v�Pca��
f]}<Z�=Z}�=����'ϩڽg2��>��P,j|���4��<�x�N�4����B���J;�*��GW�`����X6to�mx'
��?[���/��~����
��w����gm Y���V
�;����`���*�"}d��������D'�!lc�S���m�p&GѢQárM��ky�|0�F]����۞}@\ʿ��o	�ʧn�
�F��tO���7�JH�v2]���칥���X�P��MJ��Kټ���� �#8��l��!o�/�Q�w�;$�R~8q��w�L�����Ar�6��@8E\��[���J=�������>������̃B���J͖W	oq�Z�MGv�ң44�Yx����*zF�i$��ϾYj09��U0E�<F)�3�%���\�� h}( E	#V-�������g�������+3Ц�
����]����}���O�Mcw6�Xu�/.-�L�'#�ʬ����*�3��s�;,�*lк�<|Ϲ�M�$tM�R�'P���f cE(���yMDY ��-���@�c��e"� *U9��G&K�;���⯤&�YB�wT���_O�d�
r1I�c~z�!,r����Q�#����z/�/@'$i�\�!ߖ��#��ܮqF`���¥�3|F=C����E�����\N6$�@Z��+ix��j
Lk���.Dg6���9�g��UJn
{������"	�.�Uz}߹��
T6�ʬ��-�q�˷7 �=	Ԡ7��"� ��O�Jm�[�RHU�,?���W	z��_�8�S0�ɓ��By ��cLg�C!Q�4��?�Άտ��������AfScT�r�^�H����77�������}G�e��ZP���yD�_3�G�<[�t�b��u�H�4��_$p'8�E�)��P9��b�kN{��Ic޲��	��,�+�Cl����̄*�u�G��SNŋ��,�pc���L�����#������MS��Y�wض��������TA�H��W��r��o��$OɉWSտ�+���*�R�:N.������D�RJ�~?�چ�ﲕ�.�%��y&�v��_C��N��Z.�����9��8��Z�����'�4h�6��8��X�Jt=K���s�,��(�Jw/�};���V����*�z��(�1M:%�W����F*A�'���"����ڊOXA�
S�SL$o|ִ�]&��O��d�LM�P?�5/͌�ևW�V���Z�S�7���1���O.'��0H`}�ҳ^����N@oJiMO��>	�1F���H��5�vШ�#P
��&<|��
+R3ڲ�a�s�������t��"� ή��@1׫�����?;I�RE|+ɯb�V��ûɇ_5��+�@����*t�@*1�ВYz���梶M�g���j�s�zN�����}ykj�O���i�s��n��,��3\����4����e
�t�Y��,�[�Jֳ�P��9�����-�G|ػ��@L�$$h@���`�-�@��"���N��%C��8/��AΗ�����G�x�o���-�q�붳5j1��A'0S��i����i�[z���D��G�N�pG�U�k�d��:��� �'|w��|  t����A��� ���1ʾbD��߄LU�<���2�s��ɪY���!X%�:v���P�bjZB�x��R���Zy�N�F��nlG,+P-8DEO�%��+1����u����}�9}1��n^����@,�2�B:�؈j�����籣`i��� T�:�)r�젋p���=�y���꺓���7sW7�s{�|)�uq.,�ݎ �D���K��ӫQGÇٵʢ�ߡ�DNU
�I��}��Ɣ��m?�D�"��"ے�:���^7f�Tq�-q�(BfS����C�l\99#-J����vp9'����EW~�AM��ZZ��LDh,сc.	��۱��)��n���h"AԒA3괓�����*�R��~/M�4�S-�]2^ttا%UMdv|e�u:	��i�L�k��_H*?1��y|Ct�ud������F[��|���A�������K����#J�>�W��2���k���
�%�֫�C:�c��ݸ2����3���-ף�tl��Y�����b�����L$V㰤(~����a[���,�+@�J��N?�ILV��K�q��{�p�;�)�,'<�X����*�N��doN�K+/*��eJ-I�6�{�K��/�u���W{����$w;���~�W��H3q�f�⢯k��V`wp�b�$)ׯeMU-�;cZ�b��Z��@5�p�XYd[5�[�ՠ/��uӥ<,.w挈(���2��[Sx6m�^��2c�*$x�U?޹��T޺��CZ믛�Mb@�
	l�Us>Xxe�j�K�7�L(��m��S�H��t��&���.ٹ>�f���6�qw�m����ό��Z�a�x�hu����F����;�񁶸�<���?y�su��R��� )�3O���L��o���רX��m&O��~����4�΋��2ʸQ����W�W�������������lT���"*��C�����s�9�ͻ�E}�jǚ9ҿm�r �p�}û�>t�Ad��i��S�Nr�yc��/i� ;�{W��z&�7wA/�I���hѷԯz|��m�k�H�Z��F�$�t��Ps_h	�d~ށm�j���ѽ�00Ng�����#Bg����(?:�~@8_LB����:{|��e)1����g,��-4!�7�zC�E$���b-Ѹ5Z,D�P��μ�H���f{�MكU�D��)}aFy���`�R rMfSO1fs?�W���c�Iq�
һky&K5�0`O�O�dmZ�~��8!�ђس��0m6���x�[�Z-7q7�s_ ���X��� w5,�n�� {�^���̾�����ո�/\?����r2���M.J�� ���/vF���"LX\,�/8-��`l�uaH�n6J�����V���z�v��P�r-92�R�F~�<>l��/5��L��EΞ�� (����u`�ỷ�7��l�}h���z օ�� Pa�oۄDl�}@��0��b+2��JT���W�~Ke+��ꀅ�ޚ�6iD���E�u��^�'��
�SW�]P.����F>`�/jۑxܛ0�L��Q�wĈ�vr��5Y��k�8G;�\��D`�S��I�B�=3�����y��,Z��.��y�?;=�����[@t�6[⻏��_�Y��� J~�{q�}uŹ����Z���K�رs�Y-��qk�|�>��V?�����2Yk�-y�%�jpu��zBu`�����.�g�'�+  ��>�"����P��>��(r;_��6���x�_��p0�x?dW0�<ED��H)Dܞ��ʡ�� 9��]i��\^�x�9�����[�NN�D��e_k��ڜ�$�N�h�����,���5'סW�C�/��D�o��O���<��9�_���`�7���9�>��E�+ј>WMc�0�<�C9����v�לm{�d���֌�j��W�۫W���e#"t�9������Z���d���/m�]��_�'c�le�k�I��:B�­8��)eP�n��*���𮦪�K�cY6�^�B�`��]عz��NI_��\�E{��rz��C�ʡ����UAR{Yx�����ΡoA������V	��g׳}�����`��
U7�nA_��"ǲ	 ���ݧmӖn�\&�.�y	S��,��~�N���O%��V�|��px^���f�Y=�%�꓿z�I��n����c U�Cf_b���������Se-��]� �E���5�Ζ���ۚ%;�j���p��h�5�P������������勅���[t�?�N�-�e)�п$<�7��r(�.<�QY߾FWK�,>�&��ln�0Ep8G�daQ?��b<�Խ�՘J��������?/O.ƌ���k�����5R�h��ȳg��\wE}�qR��������WL;~���Mb��h�-*�-u )_���H�� ͨ�ކ��Vv�f<t��鵿��~T���X>��'����?����׊�S���wn4��9����zTB����ȩ��[.�Nح7c�ߙ�5�)����Z���L�-)�ߙt?�r��{;�S�A$Ф�H�����[V�St���@f����΀����x���+�;�����2�ts泊�� ���]�>e{Fb���^���4����@E���X �2��v��#3M�*�\y���4J�%/��o��b�A�d�S���R������P{���[�+k[�J��ֽ�+��F���W����|:U�.�z�8f�?]��,H���j]4fO�`��$� ע-�2u�%'��r���7	bfqa:+f�<�p�<Ȑ��ؘ����ֻ̦f�x(�[��X���r����lb��4����4ʍ��t.��P��m���{�<[O���=�@@6�um���(���4n�i�VH洯��d��� ���z�L%@=�rL,L��)��4~b[
U\�dԟ�l77�xDҽU����2���e ٪�Z���;m��B�v� v"3:�zKc�y9Ø 3dۧ�/@����I>����.(�k��@g{�����q�:���<�c�]C\�&�Fp������R���,�J2�a���Px	�m�~AU�l���R-W�+��ީ�3���+��lD�v��Kzu�a�O����"a�FQu�
&�?u�Hs(�1/�X�ߚԣ<�'�Zk���K�Qmq�A�$[�G��U.��RZq��8��Z��✾}�zQ�)�"�f:�K�vO�V���&a[FuGՏ%��=����ib���V;i�-�=�/f���G���v�:jk�Tұ�#�I�B$v��g�'8�tE9�Y�U ��7��b�G3;�o�9j4����L^��GiN�e|�;�p���S��{�C��`!����v>t�����Fr��q8�>!*��.���Mղ����q��?����#/�A?�H�Nt��ʞg�h����t������<DV��`D`����72��]AQD�gcH�D��)��䇶��\�\W'搸�o�s��Ƃa�er���r�f�f[���7h��c��	Q�..e�_�=�t��Q�J-��md�������DE�U'���'L䎄!=����L���J���&�Ód`�aQ��ёI�&����[�/RZ���Wѽi��G�z˒_��?�g��,w�^�ڈ"��m����)���1��
_@(�c-���Gq-���� ��d
V���d�X�񭘙a��ª����Fbld��P��l��C.�m  m.���4����WD�;g��g�
�:���~��{j�a� <|�z`P������$�����e�G �m���	���˓����o�d��U�G��_��Kن�����9���6\�i���J��.">r3^���t'����o}�E�v��W!^�ü�"�r��C���NP 7?aZ(�V�aX{'V8f�]��6,���H��bXXq�!No�u��^֪X {:��C
�uN�m�U�US�V�-�h�����Q���Z{�w^��� ^ݤ��%z]
@�(X�����ő�6!9�ۚ9�?:�����ym��W0��9���O:
�;�g�JfFO��Y�)�l� �
,��)`#ʄ[�U��7c�=��N�n/Ė��M^��W�/m`��4T]���[�تm,Z�I�~�b6��땜^*�����6�1�h8��O�Pe��S������ͬ	��C��v���/����a�A^v�'~H\])���P���_跪�4Ft�jʎ �ڿ�Q��f��C2�01��i��?�0�k�n�g���[F3?ߙ�����bs�LK�\�j�|"����P[��foT���ݜ�V.韓��_-�7k��i�����:s��w�)SWW>�O��︞t�XuF�q��ʽ��)[���wu3�Yx���hz�7%�gD׀�P�_�r�%h�m�_E��ȱ|�Va�*��6�~�0� iEeA�~Q�9N����p&7�z�t�mz˳����C��p�e���^�{*뺂B͘���m�� � �����Ϭ5�?���8���nL��Y9$�7��=��iT�/����\�!)���n=u�*������K��<��a����_p�2%��X�N�MqT%
�`�~P�s˅ W

p�՛�z̧L��\\�	�݀!h\�Y���l������8�1��Ȕue���	N�\���&>��s�������|���S�А�U�o<�w�0%J�q��x'y�1���<�,'�7���]S�D������S��������VLB�O^R�J��&��M�Ёu�5�Wn-öN}_&�R7�N���E�Bh��޸uZ �<V5�OR;j���J�>g�;-��(D�4"�J�x:�y1Kwi�k[��a{����7�۞դ����1L�3�"�S��YTW6��|��I_��w�/��c���ɑ�f��������?{nO���x�{C׳�\�ԛ�rb[�v�z+_Ax�wԣ�����+�%\3(ݹ>��$1oO�n�r�yu慫v|�V�. ]Wk2�_�c��]oLQl~��rj��z��z>�<��8d bMWEБAEeƶ�����9VT�}�`��˜�g�V���e��r0N)�yj�a�C���/��<3S�"�v���?�yB�^��;�U�/��EH�a�-��%�������^�������,{<"Ng>Z��O�%���v�7u_<����A)�(�ɉ1��g>_��~�3��^.�ץ� 3��=��F��h���`c�_~p	o���Qn��H�p�N���:��L��ÙZ@���r)?!�B���Î��QI:N)[�X@��{� ��)h-_>=�x���Z�(^��#����n;0�M2#@�u. �Q���]c��i�kU'�сơc�V�j7�  Ti���n��vY4@��)�+�Q���vf�ZV���0��Lo�S��u�g����݌:� �ѕ�,�0�.��L|VA������B�v- ��v>Xv�S�u�Vc�_t����R�I�vB
��R�z�H�W����;���ÖC!�<�8���K-|�|�prE�E�"?��h��� ��݄b���{	oCٌi��{�¦���_e��UiZB�����(��1)�=D>��*̕��
,X[|
#��  &&�`p�Z�R�a�������A�ހ�çI1Hd�7cX�f0�V (`~�9��<�N{r@A��t{=m�a�6���q{�RI).�N�� ��|�YZUT0v\l��lO6J��L0��_Y��:���)��j�A�|�E�[���."��U��[np�p}�d��!�=G�.� �r�iW
����~�����bT���iϯCL�.ۓ�U��B�8���y��Ѕ�[@��m���ܚ�]�����Y.�<�9��Ôp�z�?�C����ʩ�z��lI��n>�e����F0osSg�]p�Ѵqs�T!s�v,��Zؘ���������v�<�ɶ{n�f�ܖ:�`��X��|�@��[WQi�8�kӽ�ؾy^s�rHi������cA!�d8��`I�hеy�aǗ��ߗ��ڗ�
?����5�~�����
��4qj�'��*�H��1�� �rr6z.���"\�ӄ��D��h^�����$���4�b��޽?i�k����U׃���1���BHɜ���a'���@)Dd&w�X$�xI�w�\(/r:��3���)\B/)B~���;���|R�G|�.�w2� <��DGۃ��-i�H��������ӎj��@�����:�Vs�!Ə�k�����"����*0�k��D��|����ա��`� ��$ L>�ɋ��TYr��I1�g����={���Nʿ����0k���������d��s(���'*���A��(z�n�c@@��|r�1��8��5P�>�i0�zva��=l]_��J�Ne�CQ�8��[k�l onR~��t��ćc��C�}�>�P�u&��8�j�|9����6�/����LiL��*Z~[�C����o*v�a�L�e&p؟����w�������U@]f���/0P��8+�̣9�Q��^M"c�,C�P�m��O��:���U���n#J�q�ّ)K4Ҍ(2���U��G���L�:��QC�_���&}��{��E�5��4Fv�䷸9�ڼ�1旟��%h:oaWA�}�I�|�d�4�>(Z �%�����ɚ\a{b����k)P����3r0Zq$ͤW�ڥPܲ��̈ebn���A�5������}[@���oZO˞�/EB�8'D��~��������7�%\��c��pǥl��t�;��&���Q��L����n�����G*�є��}R0jZ�=��mz�	�j���^9�%MC)��^DjB��[ ��u*���HL�g����@� _�f�-���`�(��ւk�g�ͪ(���;�����aZ��K�g�Y�Ww���d(�$gդer����&�N䥪�7es0�5�������F�i����<�-��7��[]�xQ�*:x�Q*x."�\�,?>ۙ� �É�N�B 2���Ͽr���M�_��� ����}SBƈ-@U�@�K<0��$���.9B-���WUi�_����l^P~
e6�:S'h�8��"�/Aci���V��^ v�T�h�R�u���|Z/O
�](��8qy�3�J_�1�3(E���I>�
��4�Z�� ���qp�6��Odj�t�3�7p�h"�5�G�q$��^��IY��;5ε����0R��#ɣ�������L8lR�G�{dJ��� c��?���D�����PK   6��X��[*� �L /   images/e5080447-3a09-4b80-90ec-33743b39ec87.png�eX���=�� � " %�����JאJH#҂�*�!%C�
�]RJ�tHJw�<���W��~��纼��9sb��k�3�)�%n`��FCC�!%)���v��s��h��u�����5�r���<cYI�[��Q�A.՛�(�7Im��l�-_���5D���g1ymfm�ge�b����*�4�{hR�OT��m�l����ߟf^���|��&�N&�H2�HSx>t��m#�'|���~L]~���A� w�KJ0�|4�cm���rΗ�Z�	�k��b��iF�l�����u�r��TW'~��v�
Uc����&JR�~��@�3z���c����+����y�]x���%?�ם�=�b��<L���������e�߲�?���B���h�hlW��Ph+���d�������i�o����K���$S��*���|��#����n.T�����a��r.��<�9Zd���/7��tV�����y��O�Hd��p�wr�g}�>e���=���,߰�7��g��;a~�+��9�����6"Cp�q�b���J�_'�p�tr���`׏kk�M�͔r5'�����Djg�N�?8Vı E4��w⪡=�_5�>A١�1I��{�W�����(���}�a�i��4/J���)���N`�OgU;�'P�y�sB�AdJ���M���n��V��&ئ�I�.'N[�g�q\��ѶDTgF�C�O���c[j�����G�*���[�X����8��2I��O�������#�n�Rζ8���a���!�+zs[�B��QCUy��B��{�<�ܯe�~��M~�g'��TV!��N�; i<jQ��LM��G�=^C�;����e�0������謂!��ɧ�ˤ�{Hz�]��ȹV�G�䯿Vث^��"tgi�@��I��A{����0��I��ܓ���_�t�
ɿq��bv^#.�g��ŧ�0�U�֔��B��un)o��H�������h�����P�:����w�����8cy�:5��'�W-����"�7������r�~�y�6%��#rB�݀/
��Wċ_���&��z����j�~;^5���[| �gW��+\�׵���"��U��+���L�1B�D��k�����y�e^�XU���"7�F�x�%AA�E�Ȋ`�1{ެ����3��[��		cn:Ora�GV>� ٺ�Q��oll���6ۙ�"2�Pv�K:~�}$�K�l�s�c+�7��w�u��X5Ȥ�.$�Y���WG�����X�	t]���\RX�=G
���I<UB�)l5e�'{3�b�a>
6$��*V��@�VeY�7!/0LSK��U��\^P@c����U����藊9��yz��5Gߍ��m��'pS��Y]e��0�b�O.b�����*�D����pl���g�����<�b�O�^������6
�c��mq�Kv���BNꛧ6:ݨ���Y�n?��X����]�r���Zu<�i7��.�Ѡ�2��NټU��{n���V>�]���ևC�yǾ �zy��}v��	����7z�Oy��Γ��c�[P~\ܼ�O��c�-�I��,k��/G�M)����e�M`����~5��J=>zK����>��s�����]�W�!�g_:�1�ϢW�;�яZ�	��Ș͖�@�f�-(�p#M�ɻ��~�ߢ���8���|�a�	?�:u���)���{y�ŋ����6�ۿ�[̟�;�~�*��ۺ��ۺ��{�yy���@ށ��y�m&-U�I /Nt���os��[�a8�{d��u2k�8�L!u�C�����p���{=�ķ�z|��� �a5(���*�&(�/��.��6W��1c�s���XfvS�ⳍ.���>������2�w�}'��!�1%�/֊�w00�3������U����Gm�	����݋GF���ڤ+�5����Οk�V��ت6�;�I!��I�n�@)��&��Ж}�PU��K���V�ns��:/����\X��TYDJ�͢z��0�xu�-�:�7��A��ݓ5�I�OJ|�6�Np�#��3�.\q�<#�Ɖ�¡��`Ǿ��o��ZD���IPu��c�'�Qi��؏��i�J�;n��2����K�8`�wɷ���@"���?��4�7"�5�*���9�1�an@�It*�Rӏ8J7n��)����I����O��nz�lo���{E��TS��5���#he}<����������K�*�kf��y��zky^�
�Уu�܏S.l���U��S���c�͇A?���������[N��U����B2�(���I�~�N��tΖR����^�+q���?����o�r귡�p?|شRK	aͬ������}�*�`���A����=
�f~�36��f�=yq�V��tia쨀�G�1�����������b�Ɇ?������0`��H�*�r�����D_tS��|ƅۅ�J�8���k��~5����*�h�ZVM�0�g�_N���sYe~��]�D�7�,H�ܡ{!�/���ɢ����Oy��h+8Ѣ�ξ���{�����%�C�Q���
�-&Ϊw#�(���=����7}��]1{Y�b��Z��gIn��mGBbs��Q���7M�:�b�G�}.�&詌���$��Oq�㔿Ʒ�lz]@���?V)�)�ȟ>,�oX����������x��jc=���<�Ǥ/�H�����oS���7~�|���>�+�F��7�6o�����7u�\��ܢs&樻��M�܅�� ݚD;I�&�N��<��>P_s��Ωd���uwB%Lu��uv���Y栧~[YU��hL`��YtÏ��^���މ�������4�lOR�n������ʳ)�~��I���L+�7����L��3q�Z���JɅ0U��2�񾢩R�X�s�
��T�,��t�X����6�耛��,�vw�3������۷��A��6��ԗÝ��%��{�Kt{g�����ld�^��`�7�fX�۽o'���G\+�S5��7�C�b�fK����Ԋ���|����3M>����|c>+�F����7�C��Tl"�O QE$��;��c����u�>ێ?h�C�~���0���O�Z�a��Bu�T�[͉�l�l�L�%e�&:=��tV~����<�j�VsW�Q5'M}v�)�?�c{�Fdz!=��Y�9rq�5�57D'D®&�����!�<	{x[���F0-/4v��ip��$@��.P"�|���N��a��1%�������	�4�Ro��,��B�������-��	ݷ����3�>����}�Q���s�b-���������6�n��
j��FF
��'p��X�*w�".)ؕ�y��u�lq�b $JTTtM���~�I\/)���@k�Ŗ %��3�sX�;u�ʺ�/�EV��H\�~�� �w���`��1n?�eq�=h*��-���=�E�t�{o� 莳{�2�%̐}�߾$���y6�VI1�r���ɥy{z-�\�#��QcO��-���DK�T���aX�� �|����L���S�����xcX_[�B8̧��b�f�
�,hvt7/s!>�Bt������k���;U�f���k�T����� ��F���L��v"�kel�}&���Vy�[/F��U�-�\geY��}`�g�����O����JJ%-U��!�1�}�<����Ħf9|�_���>�lE6�o��H#.ծ��[t��O\��qro+�cI�9��5C���i��Oa+�������0�,Hr0��8 >�o�E��sv�\��@G��=�ٜ��ݗ*.�
4HX #�� D�x�U�{Xsc�����3�s���:O��-(]�N�\������J��n��V�����J��������T�.���/��A�,V^iX%q�����8�ǈ���m��	i8�?����2e�f8��?��E#gUǏ�q����u��\<�O���2��IJW�գ`W=�Q�5��UY2�+b�ｍjC�����\w��i+?��4�9 ��⌶�n�Fy�w��Fr��Ftj�^�Z��9�4��YV`�pw`��j*��^H3���E~��*�K�8�H`�x��ڼt�������D;� �ٚ�]9�k�V�s֖�[�rX`��F�2�e�_�d�������`���� Wg����%K�[<W�$����sk����赕S	Y���`�h��Y%�@�L]I2춝2���,ii����J��������Մ��
س6��o
��~�>m��i08*�9=���t�J�0	=G�CB9Y����<�qFeԪ�_i;����nl�8hJ�8f��Th�1�	��� ~���C�(2n�=dU�D���"�ɲ�o�܋e���X�>�0%��j��?�7 �<S�@�4�V]�;P�����������1
j�[ʚ�
��ڒ(��9FB��J�j�EN���x�E4G��l
}�V��g|���٣��E�d ���RgbYJ�khz��*Śz��	m�r;������It�Z&k�Z��g垙�Es� Z�����ac�v�r�:�����l�b��rX�ym�#{XP �W�r�q����?cح�͇�r}5-,�ZDs���r^\�&�އ�=MDk@da��������g� -�7d?�7�*0��a�jyӿ
v8���1�q�B`r�l�=��-��[�<*��B�5�Z~��{�u�f�uֿ�q��Z��z�8D���&��FL����[QZ�i�������e=d}�ީ6������<k�`�=C�����\8�9�ޛ�?[�;}�2�\���;�x��������y��U�=��.�����H��f����HkVIh��{�S�c�CF	z��+�K��>�CN\%-A*`;�6o@�����D͢'����eSۧ�jn���Acu:i�M5����sL�+���)Zgk�k`�r�<�J�����o��V
�q��%R�T)��#�کp�z���0ރ�r���צ���[EcȮa
��~��b��4f %6ۙ��o��'ߤ�t�,����z\��N.b6�Х,�4+A�6��'a0�K�,�29�&�`���Y��hE����$oc�F0��w�O�8W�_pvĒ�̊���r���3���N�}U''��z�o���(囱v u�[�ޙ���{�>�
�oδ��iq��%�FhB�>���ތ}�,r*\�̮�+pOcw�>nn�(�z�W3/��	�%��_j[�+�ztf��'$0��㱑͊����%2T����s�an�/��k��6��к�XM����v�^i�UP3�i����
,��.�^���\k����I�6���D�d���}�$C��o�6�wحV�8�_$8�ST�����}�v^ȪN����]�/��m{�H�`�`��6�t�3�w���I�#ql߾*\u^T�٫��nzI���L3�e��n�[;y�sB 3"�=}��V���dԐ��_�v2f����W�v�۵%6�c��3KprF����=]���s�I$���$��6��K���+=�k�݅G	Y�-�Ef�[)!����!w>Q�Z��m��/�44a��ȅ��+����/�"=�jN?��,�@��p޿�hŃm�禗�z!��mfP�4��N���6:]��yu6�	r�X�
�F-����5��N$���v��j�	ڶd:ͤ�4{��K��D7�sZeL����u��h��`@'$a�X5��:g�ӪJ��$�i(tA����2�j�i��@F���d�A=�jHP��=`�i�C!��Н�Wu��4�־~�9�Q/G�c�W�u�,�t�7��+A�ٖ�2���x��5������P�_�����~,nN�뭆��b��x�n}5$��I[��y�^�<:���
lh� 1sۯR�9��U��K%w8�gw����~��Y�1�����o"�\���X�N��a��a��ҷY�d
�ENb9�e���a�ߕ��-��꥖�W���o4!��⳽�f!eo1�X� �b�cH��;��9������w�.�Fz�jy2�)1$%�eϏ�����!����:���u{M4�54��_�W���m0�r	k/F����s�"�/G[�Yl��LHHg�Br���ɐ�x&e I�6e�P'�P{/]m��=���9�a�'t���	6�~�=�J\C�E��3����ꩪl�>s��g!_����2t�bS2g�NV����+i@\~��@瑴�Re%z�>�V@˫�TΛ0C�V�`öX��졨𫛔��ݹ5ŝ��n@��mf��]C�Ü ��cq��	0�&���wJ��b� ��[�;�S>g�a5�C;(nm0���2���q����-�૨��]3jU�h��%���<ܻ�-{�=���=��d�[v�	�y���"��l�q{����UF�(ϖ��BR�N����*� ԩt�I���� 
��	��V�v.t���[k1�Y�E�����J./��������L��b���)f0Z�\�/~�u'�� �іCAD�!РkЦ	��!���j�e�A�����@�kJ��Yg	.��������#�^�2���n��1�����]�n$8F88��
���D�q5niE� m��"P��A�-��]�{:�����Nǟ��e���5��P����!.���-�&1P������T���)� $L�L27<x*˿�
���F�W�>��ے;���0�1��!t�0�Rү�l'x^ 5�O9���eґD��fϦ:�g�7�=ݡ����i9�BKA�}B]=��+���ǝ�����.b?[��k/oU���#q��VCaaz�'����MZ�2`	�ݜ�����Q�{�#�1#î�<@{�4�*!�]�H���M��S�Ӝ3�C�^=�B�W�Nt;�+f)g+�<i�/	#�UvRΨ�5S/��c��9��o����֕�ae
�NB�,
vi�ז�M��z�5������T�Ū�ȧ�����쫛������Y۽�D]e(�qF{�p�����o�#x7�x�&pGm&t�9�>OP��O�p�C-�Llf��%�]=q0/�L�k�͐��o�>�U�tP��)�B������|Y��?����*3�dȓ�h �	�� ͦ��P������r3���xIE%�କ��M��+�_�%5h
��o�@��msx` �<N�s�;�O&��T�����n/��6�l������|�7����e��F���c��$���:���� �' m$��C%��:��YC�.�G__�3��� q:���y�:(��i�i����8֊L�t���
�0�:���[[[��{b���J`�u� F@�a�-"�7C���X�,e�O�L�a�8��ƨq������a0Dh �
P\[��p[��8>�v�n��gs�|D�|��#����A< ���6�t���=�p[��RN�!'�B��o�q<��������B?�lⲮ;KJF��/��6N��@rq�5�u����D鯋T�����˜����5�9��C������T�k
�e[�yǠT��^00� 4�T/VJ6�"�{�c&��̭o)��h�1�<˙�(#���-��(�A����b߶�)������>w`��
��O m���<�~ֺb��7�x+	@�D��@���`޹@��d��cS���΂�:RP��͠wW�u��s����λ lL5n�F����$j��5�bt�[�M`*�t���ח�Ue_k�N��ȇy=}$�r�P\=9��0�	�'�Ϊ���`s0]��O:|U`��!7fD֜k]H'�	}̀�W�l��cҗ%�����L^E���j��B�A��ɫ6��ͮ��w��oP���,V����	W+vIDQQ#}%���)��2��8��K��i#�C;�ؤ`�l��b�����yyy�9�Bm0��_��S��h�<j0O__�p<AM��VB��6�I��+��̤9��D��_�')�qo1�`Yt�C�Ud�Ju�������Q�[כ�C��60V�����M|[��<��%[$\��j/e�pe>"�{ͻ|n�#�7��Ai�+V2z���y�{.u�_������m&h�j� ��������R����Y� S����{���0׋T��淾�c��_���^RD��s�O�Ӕ�Q���xlW�p��4y��}��>Q�i=���oI����6�>ݻ���4�tC��$I��(4Dv�����'�}h�]ֹ������e�>)��s}u,�f"�|�*5����ц��NS��h�,R���:|���Q��C�ٴO���[���gH���ܖ�]sck͋_����'���J����􁥎�s���\�x>��Ƭ���V���8�d�d<��̼�x[��=�P<3Ev��Һ��x��$�z��Hn���K!�	��V��έ�J[���cZ����l���k�k���U����*�q EN��nG�R�%��M��Fh粛l�v����5Kx�|����w�b��u^%oDSN�V7l�'ٶK���[
��j�7�lH
.K��}�)�j�T�����%�Ϋ;��̈���g᧝r]��䙟��^���q�C<��M��Nw��5*�����(�l;��;4��J���+�������z����c/AE�)y��ɽ�B��H�ͣ�@�1 ��2��w
�wx��]R��<��e:���i�R��7��$��l�u���"�m?�k\j����(����펗^�[j��,r<�D�h97�ӄYfD�5?���]u��B�WD��Rlw�{+O����	܌�g��rv���7��S���fI�Bi�������;��"�ʲ�Clf�Sl�Cx���������ǔrH���#��Q(��z� ���Fz�s-!Δ�t�����ꈦ��O���O<ZA�����叼�*�l�� �HǍ���IP]��1������ژX:D/��]�J�b�?�O��O�-ER	��wn���H���ۨZ����w��&N𶮋���w�k}��x�/��^Y�]��G�xuZ4�z����
x6}68�yH�սG,��b[,\���BR}(쀄V>R�M� ��K���_�nS&�l����{�F�G�օ_?Gv��cw�E�?Ѵ��oF�Ofe��q'ꭐs�ե*f����L�έ�F��&��˧{/��G|����2ē%��s-L%kuEoȟ����.Y��u,�-�F���/�b��Ai	��j�*�Fu8��'��v�Q���v|���6�U�E�+$��$�L/ul������5]�cy�ꕟP�;__I���5��ݛ`Ѻ�%�:���
1����f��$�M�E�����,[�Иƞ_��*�zx�M��=���u�#��C��_� hh<D@��	�������u�,��������N>(�o���Om%v�[`KM�2�
,����Su#�Z�c�4��p3Oc���}�31�M��e|���bO�.�H���7p(��|���f���4;ͺ����'�E�2����o$��?�&ɘx'ٖ����Dv,h������#�|��9x�ȕ���ܱ~-DRp(md�e�<FL������f��C�u)�������Ӈ��|�Gw��dT��wIX�$G��o1?���� &ͨ�/	�ˏ������X���@��=B-�؅��H{XN;ag06V�ߘ6W�B�!�a�"s&�mo�Q��t4o������"_p������f��%+R���VǉF�ۥ�q;<��=R�F�Rb�����BI�C�$�{H?ho�a���CQR�7���J�%N�td2��k�3�#`��q":Y;����5�6U �7���XZ;�����=��pi�\�iԝ�;�T�����CP �����PN��a���+�}t��7
c�>C,#"��V�M����L�Ҷ��RzG� ����1�Q��b��h�e�o�EeS��.�Ts�A[Ȥs�c֗+�ǭ�4N���YhN�����qo�n��(�w��i��<�{���l�0'D����%�����#����z�SπU�h`��v	����W�oy[+F����o���/�V��)�0���f%y?�n[�2/+o�����[Yh�#n=������Ogg�U��Āxr�hۉF�ף$��mA��e���t���	����;�ALkm���L]F���'!��T�hҬ}��?Qh�R�I��н��J�C��)��L�\˚���iPic��d�n�yC����ѬD#���/�y��1�9���Z&3 ��-�沉�L�RX�.�����*�ن�Y:j���T��S��������n(�`�D��"�8�N����v��4���?�幨�UEL:�̝ eܒm.+��R���tU����kn��L�wM�������N���<y j��:���zU%^��"�M�XU���\I�$Yw��7�0w�_��r���g4��?��/��4�6$�k�-I��U��s"��T��C
"6T�[�	��7�g'��Z]|����aU���$Co�Ra@����ˎm�^�F�Q7�?=�G�vmX=X�O:6��������,%ݚ_��P/�v�����9�A�>�1�m�Fh�/cDHݺ�+����;A=��T�W�N��`�2},���;����5�A~�!�*S8���!%�Ǚ�j$<2�K��k�a#�ؤ�[7���JEݣwO�T/���Q�������/��Q����kޑ���+,>]R[r�g������⍑P=��:n(�=��sL}��ϸ��3
B7]���zw�6(!~�]��ņ���3{��{��N�h��faB;�9MDWVQɸD�I��|έ_\�@�K����.󃨎{7n�6j)N0D�S�f�V���B�V$T$ܮ҅I���@̟�M}<7��D��^x�XU4�0�҉jJ;�0�Ȁ��8��Z�W"��@�h��xS[ ����D���h�lpcᨇ�:n��x�U5�ʄ)8y�F�]`���
��R��V,�������ØEr|�b�~z�Q񥑂;�8(���xOa^��> �@m"�M�t�:Z$X�PE�T6�c^ُH���!u~���wr��q�h2�b����
-�2��R̥#^p��fu� <�K���r����(�d{��Õ"����qyT`t�����m	G���_>��~w$H��K��-�P�B��$JJ�I��Ͷ�w�}�0n��8�q�S�������
w�x��e@!D.�D�"ҏԏ��O�4�xE��g����}�����hN~H�^�Լ7�yiZ�����e ��dF��G��IJw���n���Ѹ]��j����r�����WsA&�>9�]Ȅ��>U�T�Yr����.�8f�:�$6�_�[��|���RǁW�ױ��Y
6��f���d��{�7���)I��!��zd�r�.Ld��c�ce�k�n�<��)�d���˧Ej��I$�
A�3_]�&t�GN*"�n�؏�x�������_1����ۋN"�i�?J�9{�j�`r�F2��FEO�� �i�}`�]��*�Ϲa�]�G~�qa�2����=O@
ӗ5�C�好I��-�R����@���ڲ����;?��J�N��ꂠ�l��L8��L��r!Mb��꽤l�"�}�FFYy�@V�H/���8�Rm��{I�C""	ꬫ�Z��(�=��I�e���zt ��AD4Β� 'ܥ3��B�A�:�a�!8�j/<r}ՠt>�N-���_���6��82��v>���l9c���?w�Oqs�j��E�S}z��A��xX[Oծ��J���q�=��U��*>�8ic����������Z�7B�:vS&s�:�+�ȩЪ~�7�o�[[��j�,�b�ó\	�L<��������	M��#�~ꀪ��|4~Q����:�k��\i�ws�`��D��d�i�iL��{*:"�^�_��2>t5�N,�Ȋ���vw��*�܍D���~��q�Dv�:#�h!��R?��W,�TO�C�f6z����lK�DttE�P���E��������#�}g�I=�!��%q�	����S ^jc�H7�V� a��(�v� 
���@���v�1��z�r��n���)v'���w8Y�B���'�!�g�B���_�Ѱ�I�g�&�e>�K���B]����o[����#M�4�@?��F�e�ßlRI�;��	���OF�Oi�6l{�>@	��)�r/�c��>d<yr@}��������K����<8�#܏2��D̹�!+�x́��k�'TeŦŵ�:�d&����bs�����C�H�C�g����"�`I�ʈ�1vӗ�ҕ+U�*�6޳W\�{��lg�߼�ia�8~����2��P�iMNJ~�p���)��!�u�O�0{��e"����fP+%��HE {b���,K�~�*C2օ	-�B�n����wQZ?,M}��JH��Ct8��Ib���!@�~�/�L��}�Ia����%
i��1��p�q(l��X��Jm���������I#}�AAdqϢK�B2�-SO����'>
�(_�Ze���;Aָ�S�D7�r��%�c�3��)"���s��7n4���HF��}�ɢr��/7F�=>� ��۹"����V5R���F�@`Ok�Ȟ� �ƀx*z'��*�W&2|/�E�a�*�#	�w�S���}�=�M'.ª'/�K�0�f��5��$����s��D~���֪G�ω�&B�w(���!��5���f�I+s�Q@wo's:��&鷐;[�A8�@�SM}����X�	���Xa�z������tP"$"�ҷ-��J3K��?GG�ɋe��9ô"�6Ǔ0��?=�����Lm+yؼ�6�y7�Z���U�������NI���/��q��o�S�k��ѭ%�K:a��i'��,��sfSW�G5�,�"��H@F�_�8�Z,= |�3��mn�d���	��e���,�� K�E�ejW  -��	A���+�	�w1���uG�����o_3���v4�?��P͝h��5_�
����h,�D�n���x@��;j��4ǣA�e��uB�������n^�ѯjˌ�m��+=K�p�����R�;�8�,q���7,���GNO0ܬtɿ���h܏�e-%�T��B<�r�x*� @��lsG;�M�wn�-s���N����s���Ze=��%�Q>=��ڿ����cZ�!|a��Ɩ����{-�0q��,�m��@<vW���x�����E�y��:��aly`����]��uT��,eGȾf֯>�����p�9�a�����δ`�|Eǅ��g�������&��&g{bs�PV�,2�u��t�bPZ:M�\���k�m+����m11�m��E���h!�h��i�u�@������
��e�0�#�b�u�\�j*�>zG�����/��M"2sE�@�Wo�z,��F<�W�y}��6Т����N���փl0�MBM٤AA�x䵗Jϓ�T�]��5�T�\�~���Iw�Q��淐�ox���6����O�I{9���Wr�ч�n��X�����UD�m�KR�w�C�Ot�(�#n��oXE���<�waM��u�p�p��K*��h[,��KI�ӗ*��nhD�F�������yUG=�
:�#�R">Y%��O�T�7Y]����2`3b�clPߒ���Mk2��N�X��@��$x1��s�Ƈ���㈋��"��r�|����/nL��`�-���߽� �x�����f�7 ڽ�QB�U&uw�k�+H]q�.��Һ���Nt�L`9�	99�F+���(�uο-�⏊�ǩw�"m��$�������蟸��CmM%)�ۻ�+n���*;�C2z�%xgo,8�D;����S/MH����{*.-��D���JQc�j����_��gD�8����H�6XH��v�ʉ���ֵ�B[�KezE4�֮�5A��[�F6X@
�\�|�"�"F2�j�vv.������̮��=-m+K��M��+��2"��X��vS};mIsW�F[��ڂ�a�o��ފ�(�Sm���Z�Q�Y6������[�+��q'���]���P� �ԊOK�ފN�@�/. ӟ$�|8��|�9��L����~�s�y
@���đ��r?�鏶y�<��f���^w�Ft�ƀ:�����Yk���G�=�����XL����W.�OS�5��Ɣ+���y����$�
��v�z�SL~���-us�s���*J윯��C ��]E��AN��7��Ѥq�9�~"��(B_u�7%����?�I�3��f���8K�"U*=��i�n��G2���u�K	?�BH
���u��G���u�2|)�Q�u�V>.��[KG���c`��j=d�C��4փ!��iʾH
�z��Xb�_/�H��$N��V��9�������z^+���4�a��1��6���v���*��[XF�t���W��Ͻ+��&��x���U�_
�b~7�?q�<��iԬog�*��n�=�|�0���)ۈμ�,��?e��<� ڱ��XֆFQ �:~Y}��\�NP���e��q޾^g�Ԅ-�e�%j��K��>O�a����܎D]��1�3��z�u��s����Bz�H�C�:��h?NJ�<�.�ײ!ỲR�9,�^V�ˊ�(��ٲ' ���u\
O.n�`P��������=��,撣�V+�o�0�*�H��B,��5I�{����F]��}��֖u��)XR���B�vǳn?�7���el�ʸ�o�ɔ�^�܅��+�&3xuۻ��h�p*�D7�wp\�y��^,��?4D����t��%�%�:��_&M�:�7�:���i�=�V ;��aT�������9a��3�X��J]��joD�!N@<JC��7g��Sb-�ܸ���@=�c�]|�Fd�<���C۫���>c�n�N���Te_�r�5Ɇ	�q�C���p}����]k�5��bB`{�GŤT�8��#��*���M��^�iv�N�ok,~����"�d,��v�A��l�ޠ$�{�SP�~��&����X��� 9�Y{u�Ji��7��xG0S<���h��ӟ9�얥z����	OO�,\nK��}�9S>�`�	+�T��t��x>]�ݩkѐK�@�3� �A���%���A�!�K���2px}\�H�� Ks���"|�eb9�*�k�>��2е�xო&�@]��/?뺻aegW����=@���(���X��A��4' ܑ	����3�>�B��4���Q����q�d�y�-ļuSY��(��{�л��6ҽ�B�*8.˼��IB��*�^{BM�G6"]k����>f����4t��O`A��J�~@�zXy�[���|�X�ˊ?����il�9�ż���Ӷl�˾O ������]z�6�8�/_��Յ��KL5 �.��ܛ���|���'�)����q�����,�P#�@S���u
�~0H� %N#F���B���Ys��c���'�kM��e��>��8� X�RF��YY�%v>6gۖ�/�1���^��}�QD5~mv��/Y�x�C�@���y��ǫWz?>Q�?Wz��QMl�)!�3_�iQ8�m��`��60B�}�[�!� '��#�r�>�Y%sK�3�N��=�J���������αr�({���U�gz-���@�����ɍ��X]�|Q�vw~|F��2�s������뫢��ۤ�$�ʽ����E^�Nv쑟'�y�6�gO�c��/P�nx���GO0�c+//)0?�Vj�M(�u��d`�oR\;��!K��������ٍ��-�*)�0�+�j��rgʊ����6��)&��q�l醒F7�0����렖���&B��Q�U\y �W-���m;��Dg�%��*%�(y�0�:]��y�����+I���ю���f&:0�v��-̱H�gZ���Ke'P���\����N!���u@�>/�}�qb��t�2�!��.�Ѓ/)��m#�2�=�ne1|�p�t�Sy\��!3���K��)]߭4�ݞ�V<H�@�?����M��T_����mD���%I`�S��M.�� Ϳ���cY-5���x���G���qqcl�f-�z�RN�D���h#޶�4&	�g���ч��D�o����jY	��/��!�>�>��|@�&�V�q��c�]�{���`X㛩v�,Եd Xڢ����܈E�`J�y�}�{��J1U}�̔�8��рT'�/[e�R��bJw}�r";|! D�$z2��ü�nfjaVl�q�P�Up�"d��Ļ#
�,�����XbA��Tl�i}m����c��e���X����m��Y�=JA����7!��e����!9��4y�_�fj��O%wFڈk.��"W����'�h���L�%t�.��𓭇���$�Y*�0��=�#7����}�rYZwuO�$<<�Db���M�dCݾ��SEn�BM{��K^�F�>�>��&��IgD"��K�\��7E��&��#���'[=b��(�$����Du�{&��^��9�hy�
�מ n�y5�E!H�P��}b	�=�}�-ۂ�~k��^���?�n�1��k�c�=2M���	2��!��a�{ԗ��!ߏ(%��%3l&�&����q�>/R���l�A<�7%�| 
���"�4�Y{�P9i�X�Y�A\�t��i�m40)���q��'�HU.��j�cs��vd��{�=��,��]+�R�w������"VoY,\A�~֜�(M��%��d8ͼO�O�	�U3l�W?u�+�7�����'�ܖ�9��&�5o����,ɂ�ki�0�_��na���A�>	�������@N_₹��ɮ���l	�	�f~���S)M����A%B��|z������ @e<ͦa��o��1I܌����"D7a�WD��f)G��2���������:�?R�Y��t����*�Ǽ$s�C'�e�V�Gf�r�_�������t�%jQ���'y�1Z��Fj��{�>5�!�N_��-:n��[2O�O���׋t/6n�]��~��� ��w�㎧�C>�@Ot{JHˌ��C�*T�,��r����2�_^���<�ˑ#K%�e���QF����
���s��Ρ��v���@�-��w$�����}F�vj�\[�O��<��?��J5|]����.�bM���Re�!>ȪE��~��F=D`V'��D��#?}�f}ڔ���u��Ÿֵ+ ����Qޭ ^�2�L�^�D�=�w`m�Ok|墖;[l�q�o��-+�����9=2��N���n��{p����x�?Z�f��ӱ0uD�̝���UlzU�٤�k�4R��ߘeY��w��m0*
C�/?_��^nLW�D��ߟ��h{�����ԏ/���{���j����v���� �UB1X�r��;�����fe(��-?��¾>|�?�;~0�^�Q��W����R�2��zd���ꡛB��`��f��ťo;_��|��Ȍ�
6y����(À��H~�
	�����|,�*7#��mAD�F��?�Ѥq<���6�^@  ������ʰ(��o�PR��0�p�.i%E��s���X	%���Z��A:������������=3�|�̙Y��c�qq@h�`�y�Bs���3�dpF]i�ǟR�}Y��X?O�̘m��49���h8u[�V�x�O�!�Q^�^Fώ�XemI��,ߨ�!�lVe8�j���y7۾���ꬲ�l�嵧>�C��(���5��W��TT�#4��+������HE�(���$`�lE��¼�q'��4��2ɛ>�µ{[ �1�� NO�f�X9�The&�1dϜpH��������j�2:�����'L7����O$�H0�RX҄����1y�<��,�/*ɏ��&9�n�j���!��h(+7w��j~u�|nѻ��2�-I�ﾼc��O�Wl�����;�`���Ԕ> ��͸s���w��F��ҫr��i�[��E>9`���g>�l@*�x������p�{��.�OI0�|1��<���~J��o�^ȰP{�*F����͸y��_4*�a?�i��kb@�56�Q}؂"R&]ҳ�x�����iGT[���:�uP��c�U��Z+�۵X՛�����hL�m�� �t\�M%��_���+&�ޯޫmxػ1�lf�6ʫ�O��W�,\�ȏ����Ӄ�ގ]���tD	�ڷ�E��~��Oә9y,�9���k+�"���/ɜﴚ/�ʍ�9s��й=�a�T���Va7f�8F��B�Җ�ԗ�nꈁ
O��؈��V��~9cDq.�]��u���X����X�m�+Ҵ=���s�~�g��f�0���'hA|�>���������0���^��Qf�W0<y�S
fd�U����`��n��83c&39�y̍Aβ,%��Gً]z�/L6嘭$� ���ȝ-}|^�6ű��|ӄS[ಢr�����@ft��Ovڜ"idr�j���wU�o��ƺ�6.�<_,�&�`(�F��q*
�ò�n�C�WP�x�Kއg�@g�x��P��mօrW��8���_��޾N�&���jz��	�y�m���^@z�w�������'��&�Y?-��KP�
����o~?X7�ӡi��F��s�/���ʺ��
�G}�=���8`�
��g��B�W9��M�j���P0KeE�7�ï��M��9D	�X�y��j��5~;�es3��#���F�.(L\g���yk���ֽ����l�c'���>�S[�wj�F�vb� ܍L �=0����Զ5�?t�J��׸;�+���Xj��M�"+1r�O��3d)٪ϫ�.*󺖳ᵦ$l��X�BI�κ�n���~P����wߒݒIU�-��[B��j6V�m�D*�x�ߏ"R��s�Z��?c�O�M�)C-շ�퍵5Y9'9>8=��R����*+Pn���G9�(�I��$���ۭ��A	�	�T9���x& ��tRx$>)%�����/&pE(
�����ʠT�[=�_����cc>h�1�FS#Qw `-��*����93�)�N_��k#�Ha	'E��_��H���\��S�@E�O�"���x�y�����.b�!�a�ۇd���R�=���>�cV�2)�~J�G�)��[<얨�����en�]SƉ���ɵ{f��z��YǏfR��$>m���h�"M�Հ�J�w9��}d#�ƀP����㣑�Y�Qs�%�!l4~�0ԠIp��%�ג�;�Uڏ����n�H�i�������E�i���{�Dfo�>$@��c��C������L�e��sN�])�?&�d{�����W��0R^z�֬����5������F�\vz�9T6������~�� ��oݧ���|��ϳ���O�Ml�8�o6������B8mkYP�Y|_���.YEm��������hP;�*��~P����\�ln��$F��4���00e,;����P���M�=����;�X����o<@���B����8��r�s} /f-����A$�����e/����
����y�� C�.d�Fglb�����k���8���c_�>�:�mh>k�� �AI�p�P�:`��l���㧡yIq�`�����>��(R>��p"��X:�^����j�`,ƻ�:�!�xP�H�Z���s+i�vUhmԸ����_g9�L�>���f(�6��C��)q�NO�	3������Tq��s�bu-p>��~��EG��'T� |�sN�O�vǹE��o�]�y�d�`�����,V������
�e�Ru�����C@&>)�CW�
����K	�5w��q È盧Qq��q���T�ΐ�Ɇ1Xt2s}?샄�|x�ǵ��1�i�i�~�C�͕��Gݸ�ܵr��.����q۹l� �E���S2o�q��d�EA�[m	Jϱ����G|���(��oP~i��`@�X=�جj�R�N$Hˀ��z��F`�e�F���0��^���L�Cc_g���v"����������HZ� 륩��0eu�����94���л"�n1�i��7��<�ȭ}��bf{���@�!��?*�*Qۯ�C���~5ol����ς�*�j�b����+����[��'�ੵ� ���X�����F;q��׷'��_y��p��6�@Eš�8���~��u9l�-�8��>qKEgh����P-XF��eL��)��\���&/�����{}��ؿ_�ڐ�oG�P̱h4�+���-�x��������E_�͞KA���?�=��@��\���3hM���f�	�0���v�t���|A�M�G����c�5���i���1wY�
��l5�Ha��i9���r��p6���v ���7��C��M��J�cH�c ��}eGd]!�G$�56�R�@���ڲN?)�Dpk�mq��Ȯ� n^}��"����� �_:�J��t���"m�f�����k6{���Z'�L������R�fU>e�w���+�T����X/�*�����M�h6mCcP�,�P֖2	�' ��7�S���U#Ҏj�"�
R;����()�ee���0�I�6ON²�l���Z[=7#�"͠�'�Fnh���F��� ^�|��|��@Z�������n��������Е웂�O`<��:2��'ό�f:�J�����2��9�X|�;Vbڰj��S�v��M2��.O�z��?ғ�WSb	�dP/�Y��b�RɼXEc�E~��g&)?~�to�S>��O��;��w2/��Ѽ�3M\�Z�6mc��\�	YAS���ɏ��}N�w��C?�s0�������N�A܈@i�P&�Ւ��%.�f���
E(�㦵+�ţDV[�B0�W�>N������aMW*�
�Wx�Ld�d�سvnɼ"����"L�]a;뎪|�γ���N~�\�1~J�z�ǖu:�Ǎ���P�/�p�S��H�Rx����1��&��xӷ�%�˘�8L�! m��j��͝uu^Ҿ��U9��z��>-���7���3��+�{
]C�{�p����f�RZ���x0K��o�|��$��{�$K�x�ԅ.ÂР�8�[e$�GW��I�b��t���l��G��ǳ	�w��{Ku��$E{�;������K�W5�dgΙ�KO��BSn>�[��v��
Z|�4x���%(���<e�{J��)D�3%J��l$�Y�c�"��[?k�b`��/:��RX�`�~�E:q�?0%�}r���QQ���A�?�k��&���4L���$�!x��E�FIh)�To�s4���ui�Za�,	�����.*GC|�u�U(A��U8業�n��܁�M��s��W�د����(���S�c݌i)����'��ï���_K�	�ղ��F��0�v^/꼐�X���6읻��^ď=�,���������7~����������LO�����+�I*���b+j>>���S'3G��V��l����,�%�Xυ �s��@�^A%�}�d�}J,��Ǆ���)��S�M#�%n��l�-@�y<�� ��h��2j'��~��<��G3������Y���w��D� IA�}���bn:��V�U3�W�\�O��m9�-�ˉY̙�	�����sw�kr3X��a�o)E��f���¥�"��E�S���+ò;�1����3���*�����d��������,�pI�mB-�?���r>�S���R��O��!����A[�����)�-�"��DrN�'��j����eۼ�c#�i��:ct�;`R�Y�Q�9\hh@ N�zj����ot�����۞H�h)խ��h<ׂ�|�y*
�CS��!��ʧ�\���k~��жX�]����q�U�d�x3_�@u�_��A�@唱t�`�C���i
2�����TNt3�ܴd��G
��������
�-{�-?�ԙ�;�1Dc��9�!�QN�K��+��J.��t��;��x�:8V�Z�A;�aQ&'�	�[����*���2�lsb%�O�/n�J X���X�e2t�%�K��1�Vl���e��)�^�@W�&��?>����zj�7�!��&VѬ�h:���
�h9;��A��(k-��1�L�++���G3tI��Lu?��N��$�"*Cq���`����F0s�@������*o�'u���rH�z*l���gE�0��\oo�`����j��4�������b�~�c��<�Rm �̎�ף�+�3J��/�93����}��dɖ�c�_(MªnW6�1 [)�@�"j��ґ!�([X&���^Y� ��d��v֚Yw@���i�h:7����P8h^�H��j���d�L�����ջ���N��Y_��\��c�n�2K�B0��KBt�2_\ӿ�A�Q�l��	q���g������}Ew̢��I�i���Y�p��׍Z��&Y�o��]�K���F9cez�����tn����q�A��2�P�z�ӲD����7)>&�)��o�+�ft�c�k� ����.�a��u|4�X�Sr�Z��WisH�<'8�~v:�WOTO2���
;�M�S,G���N�����敦/[�<���n@88����(���*�J�<&�� ��:f��ݥ�.�H~F\����xSpv? �X�����鈉ᖉ��Sb����|��/�_^PC�4*#�n9N���n`�r���<i�l�	K/�/)�x���=�;�e����R��k9f	?����z��/��ٗƶ�E�{z����>r]�H���<V����?jk�.���K*��+WlH�؃	��M��s�<	��?��UOp�&���s���x������LW�o��m�����k�Y�w����X.�#�$����K�'���:{ �@&�I����^Faҹňl\:�;+֙�ƺ�k�8>#���,��a�XZ�	��o�ys�^$�0k�v��}�"-Z��,!l7�
���7��YN��)��!�)�������F��\_��9�il�I��j�X����:nh��o�r9�g�0m��ꃺ&F}t�f#��H7��x*���6���`b�t�q��3�Q;Hj�չ��{�|��� �O�{"�D8˲�e`�hD΋++���'83�z��ˣ�J�t(Ge������7>C��-H(6QS��y��������?��Ԧ�ǩVLQi�@=�(���O�(�~S�y%�4�f����U�e��_�j�����l��\�ZG�Jش�N�w�K~�irF۽l�9��{]a���L���r�y:��9A�"������a�M����"����y05&��'	�a��s���y�[�1ƌ$��R��Z5Y4�A�3�=�*	D������!��=�z��ɜ�7S�v��gjK���2
1���Lh{,+��u��-��0׷Ig��Cҝ��N��y��\��3�?���6�|<��2��}��5	��b(P_�B*ɏ��ĕ�|���^c��@Tj�0�lXjݯ��j�QM��Ï�n5�;����XU��$�D�D�P�b�sǢ��?�	��"�}�&*x�V�⼧�#�V�����TB�Y���P�ɢǤ��C���2�o%�(^%j���_�c����\��'l�)9�.�I�2?n/�O|a7n�B�z��P+��fz��?�l��V�*�jj���R�t�
�f�n	�5붃�����t���|eEQ��lRr������:���$�MA��P�Cߝ������'d�/��N�{�����̵�K���YIH_�b��ǚ?B��y�	��;yF@�C��@�d{'�R~m���o���wr���?=7A�b-V-#�����.�j.�Ϯ�0�ບ����|����b�m팲�5��}�'!�
�v��2��¥���w�%��[k5a�0]�pҶ��.��aDFUa������Jᐌ&������{����V\d��L�W�����a���/�ݍ:���k��#�w�4|ڸi]T׏Cax�0@<�
�b���ሁvHC6u<g6�Zm�7�)�h�L�w���ӗN��7S�x�����-�� ���?��Ew��Y��[�~3�tA��DI�BB�f峰} �l��d�{/J���S,'�� ��C�T���uL������7����N3��I?f/w>_u��,t)ԟ��P{�:���/dY�{������,T�&5��&)��g�ݩ�d�vmr�*E�Mկ���yEmg�Z�h��t�%����	�&+k�p���]}uߍ3�����4��}�"�A�ZIWg�d�?��-r	��h�2�>�����ἦ�y�u����[|�wB_-)J�����~͞B�cV����6Rv7�Wv;��{����E��14���h"Yc����ݘyD�H��>��=�6�t�����q!H꺦�Xlk.��U*ӥ�B}��7�;$���; ��;�ԭ�8�n�&"�A���
G���_�}[9_⧲���X���}+i�:��+���yd�~��n��jﰒ)E)���\�9~k�:}�쌙��:4;F��117�!㾠�	���5�d�^p���tw��_>*�;=�il�Y��JM�hEz\�ʬ[�~��MȠ�>=�;��]5�.���<�͞4�Vt�*�O�<c|��>�7Z��e슨~��x��D���n�}�\�]��$��O-��OpZ"�x4=�À5�u�}C�:�ň���祭��H��~�JuA�vi�z��E�r��A��B�F��zk�=烁���9�k����09�c�p]8[����Tp��f
����k$\^k�(�PE����,3U�}�1�X;��I�_����P^�~�]�b�rp�au�-������o����*w��&#����σ����Vǲ�`�>-������Pk��E���ri")X�T�D%���F	'S��8�`Z�v�����?��q�<�Ѩ��o݆�dr@	R�[%��2���`w�|��O�]�c�b�h�_��%�J�
�)t:mV����;	���
S2p��T�f�}�x�-��͓t;��r�����Z�ķv�2Q�/e^�T�ㅍw�H^�+��3��VM��9��S���L~���Q��7B.�)�%a6)��h����P�hF?�� ssz"��̛Q=�r�$h�� ��dj�F !N�X��tW���)�cRق���
�2ti��!Շ�MbW������h����KI��s)x�;�����7@�����&I�
���=v��4�W��D�$p!E'/G@B(b�36b��_���v:p�W@x�3�g����"�F�7�1ڣ���MC�D7y%�?<a�R�9W�-� ��t�t��fZ�!���#�ҫ���m�p�a~U�`�x2T�/���C�.o��w_j��M�JV��ܮxm�)ˌ&�5�:��z&�r�����O�x϶�"<��n��y���}����t�}����!��~���QS>J�!:�M|!iU.�JUcH4��{wu��:;�����*��Mӥ���@��u�jF\,0�����}lȅ�j�֡��w��C󓾝ۡ���BE�,\���[�K&[Sds�x�x��1���J����%��#��Ⅻ�8{@��7~vNU\�<cFV�_��ɗt;ӷ��`�	���!�P�)��r�]Ma��<�7g����c��@&
�yb|yÊ���@zr��Ի�~M&ԛ���|<4j�I�	�.��ׯ���Kc��A6CW�����Q����_&:|R�Ϥk��o9�x]�)��c��4�S�e7����4Ɩ);B�s�^���S�4�֚!�����hb�O��	n4���K���c�\wD6my��>���k16u� F>q]�K@=�w#�e?T��iR���G�s��p��PJFֲ��#mNRЯ���B��UO�,D׀d���/_�O�	�|�%-�����܈/�� �z��T �� Z�j�*��|Ğ2s�����Uը3��["pͫ�M���H޿���5'�\��Gp�h6O�u+��_�N�ܡ�9j:]Ua6��G�V����F�����T9����~�3������#�ߥ�-�4�<�o���O�T�	\By~K�+x�=�Ӧ��<S���C�še�N�b/;��G���A�z�(���<j#��x^�ކ�h.5�HF��z��(�״���=��xg$6��TȄ2��v9�zs��:֨
�-ZBU�X~��m���X�=ݺ��� ���7{���P*�Ns5�Ww)�U�2���p��f�H\c�OK���|���8Wcoa�\��.�A�kU"~��=tī�5a8�W�ݑ��-ϵ�ү���Z�_�%S�<����!?`�M+턾|�g5�>_�}����uB��9i8`���h���ؽ9�
�N�V�(�{���0�/���jz�`ڏ����E�3ځA櫏yw�b�o���tsx9�RfX�O^'^�f��1�����o>w�gY���3Y�ly5:�)z}Ox�%�N�`�+�J�����g�;�,<�p��Z�D��Y?��^����t�H�V�)sf��q�VYC$*7]�T���&�Z@�+�eZՍ�����:�B%g]����(��?kW���O�I�=(��;�7�e%DS�\�Ζ��i�=�Ejo
�Io�]������qRk����CkͥF}����(�����J+�9/W����NwEr�Oxo���);�ṿ~h�mD�}�qVWO�Ǩ�`�c�%E���gv���A��ಁ�]�_�e�־򞌐0.��!��/���4�/����P*�۾ֱ�h��3Tz�:ڛ��.�#��Lco�o��t.a�Yʏ���h�4Ǌ��q*���ړlbΒ��W�_��_o�h���_B^��1�t��'W�D�ϐs��[�������ȰE:tK��jQ��U�'7~�#��L�����أT�{~��%�fV �H�󄱟��/�{l��r�0�?��F`cU6��Xf310�B9�X���u���� T������Vp�
M�x�۬��bo7y@^ƾX8x|�W2��j_���3�~�p]�|�ꆍ�Φ��ꈹ�wH���)NK$��6�{�գ���osH��vJ��t=�w��y�D�V��v�q(I��n؏�I;���S�$�c��+g��oߢ�3��&��FB~$�һ�B�)��+��h߅�mn�����ǟ'|a��(
R�	g��[��) g_ʩ��*.<gv��!������4��t(��_}(���u"O���
�w@+�ٍ�2$_\����<p^UK-��Х���WB]Б`ݕv� �(�_t�����Ebޏ�]�ލ�/
����@ᠡ��!|��<$��m��5[�׼�!DQ��s�iB?�Zr��w�����J_���v��}=��4�ފ��oZ�X0{#)�X���dp��w6�*��dcd��`�~x�O��/?��W)WF��S�ݿk��Z�#�,;��q���P��զ���y�O��ĂY/pCx4��!/�UB�������~��-����u�>�E�t����0� 8�RA�V�[������5��!F�<�K�U��(�0�,C�h;/��� ��
U�2�ؗ���Buq`���r�t���8⯥5/$��4,��m�Ik�y�1�1���J�9�����˹r��Y�&丌��)@C�F����C���L���m�:]�>A�"@:*?��K�5`�A �Z,�l�G��;����Q��N-���w?��tW��l� ��}wu&��pdU���t��5����c�[�:�fK�'t���T�lDF�s�h�ZH�{�I��<�¾�24��-_�o((��ud,s�|*�]nMǨ�[�\��B��)�30�����0nO��Hg2[F��;��f�z=�>���S�/�+�h���B`�`z�%�����]�-���2�37���3��Y(��T l�/�1E��c����c�(�����ƤWe�D�}�U�G-���Z?�ļ��f^�C$��(;G�s��s����0D�/C��ݮ�`�y�c��v�jm�k��^&۝���vN��z�x�����ԽU���e���x�^�;�'F��Z��J���b㭉�Z?�������U��H�4
�=D� ��</���G��4գSM0�7P�?	.�<�Pٻ�#����T}�F��)� h��9]��Wv��0���c��xz��l��ƄR-�<5�֌hf����e��Ѥ����|����� ���+�aq�x��E���Z  �I����"wb�F�g����5���i=���Q�}��}E!��k7\B��̢[)�6�ʊ(��z�W��O'�s���?Y!~s��ľ�TK6��+��`�V�t: ���V�\.KJ��b�Uc�[w!u��4q������jZ�VT����<Z�NA;�wM���`�3��˳O���/�5�0����L��rLʦ�Q���f�"3�'�_���E"B�I�a���sm��u{ON�(z�=��<�4n�ߞ#O�Lo��4t;i��[&�� ���o�(D�m������ɲ�	%��# ��12D;t^���Z�X�nSY[�U��2B�P�,O��iŀ�OP���`:݅b�����P���Y��&
���[~��#B~�LڋL��p��M�������|f��zh}�G]�1Gn�6�uW��k�n+�q}���?�v�.��J�c:_F�k�u�)�]�32�$�SN��d׽F?޷j���A���������z
�L�;���2�}�)�Ӳd��ثI�i��',�sԺ:O^�b��nyw6w�AU��I�@�Y��m���\��[ ��06E�#` cx�su5�Vx�DRQ��zŎ�:&�FJ<NU���`y.x����B�����:w!��l�p���ߟ2�!n]�>ש��q!�|)��P|�����o �u�PO+�b�t�+ML1�0�R��7�Wo.�c-��
(���������R�V3j��D�{�&`]bj�ZY)���������CUj��z�ݮį��Y�W{���&��&R����U;i�__ݕ׉��?9p�?Ӏ��27e�1`i:�/��2hN�7櫞�j�n������9�0��-ٳ�Z .�@��GE` �篺	@�����J�%���`����κ����Iֳ	(#t춎��A����E!��u�8�ؒ�nr;��OY��_���gҷn����)��!�� ���o�zZH��n4�#�A�.��������?�����[Xa	��O����1ϛ���~��<���J�*�9���o�3�R�/$���*�>cp�׵�W�w��K�#��AlA��U�A�ܷ¸~>1�s(9S��C��L������k����<�U�KB��$vmy��$L@ie@0���wB�_�۪(���x�1�Cw��a�W����;_HA�pnzpcI�߽����Q#�K�ka�kQkQN����$�ռY�d7�� <��_�RG�\s�Z��u���^<~$�}�6뢶$�+�h��"+23._ϝXx�#'Eu(ϱ���)�*w��u�ó�ErRm��1%R�|/*&�N/>���{�Z��0�{#�����'�#�i���C�m9��<�(Ě��O�@�,�C-G�
��jUlI����tb��fzl��dVV
�*��dL�/I�qNi���,����W��G	,�<\�N���=2�_��Q�����a|4��(@��r+�9�=^�ys�v+W?`Ӱ^oAwD�iX���M*B��������i���O.����Q�I(�%F�i�Eh؏ X^���ą*� A2}��F��d��$�2����;���A�����ހ�&Lg���y�|=,��� ��@L?e�'���wI5u�};=��B��е4�g@���P^���5�⺰�:K�n��j�'�������x�m����	�(�?P�T�d�U�{s��W���U������M�fo�!�p0�p�:}�,�>o���FI��\�?f)���C��[km͕����Q�����rQt-��:����L�
��%oO���(�#ҀF��r�B�W��/�Nu�����W/2<�-��F-	xF�ؖ�hඨM��O^��`b����Z�-ʢw�=Z�3�[�r�*c+m��(,2лvsÞޞS��n����O�;M͹L{:id�'��'��@4Z'(�Y<�}����4$�H����U�.�XV&}76��:e�q�9\�����Q_i���W���Y����֣R�D��� ����!2�x9O�ގC~�in�p{�4�K��x/�.�$n�r*�?	0�� ���,����+����g�ll�b2RDX�9h+ch�i��+�?�Ȓ�5�Vn;����	��� �&�0|[̇Mqb� s�$����p=T����d-�q��a�TZ�����iM0���AB�|�G�p��S�k��?��A�nh�ߓ�m�L��ĞZ$����,Hf���<�ш�=3���G����^V�HO-(ꥭz�^�c*k��0�������##����W}�Ǐ��|��~��〴{���wD�
���ˤ�A
+���~�w})6��{4���$2��+��H�E?��U��������];7�G4�߹�U���Q�lD��q�����~c`���`⬖)OEx=}���r9�V���ߟa��+`q�0,�[��]ɶT˹(Vҍ����u\Sz�jZ߯������Qq����
�`K�@�I�f7��K��y����F��Ib��6#���\�\��
ᴐ�\��(�ŀ��������W�꽊��@u� ��*I�qz�Z
b���rx�0�{p�g�k����Y�l��hm�R�]qؾ� ո��^B*�L0@�&��ķ��E����R���|����mN�Bؙ�$_s G�a1�+�on�?���:�*��Jb��U��mH㴚!wR0ܝ������YN��0*�a�EzHb��|��+�ܪ�D�
u��X� _`���'��{��Wެ��~����>.�C?�8�j�� ����V'Ӎ��>q��n��)�,2�i�tZ����zp���i�4 �L+-�E�N�K�=C==�C���[������ү����?6���|�]�:Ϛ����@�@��|"�:c�}Sy��ԗΌ�� �apg"|H������T B�3'��,�dQLc�;���!:���� ꥄ�c������H�����S�y�wS��O	 w�������]�˹4�Qcr�^\��,�^H8l�#3�"u��j�S����������F+��9���L�)�s�c��D��t����?��Q�A;��KPo��٪���(̤h#꛰G��甸��̫)�hͻZe@� c�֔7�K���@w��׆�~�(����+��k�]|�n�4�%��g�� ����x�d=6�*�ɽ!�\�c�m-F�&S�����.÷��Q�G�����w���o�'t�da�&��`���)��
�C��q����)�0�������_�!���n�ւDzHmـ'��B��xN�ʳ�,�Ԙt���f�#?�m8d7mD��g��[5�P[}&���ټ�h���}9�JK��ոγ��CW������-���&>��\� dg���<%l�<D7',S������e�1Nq�fi�p��J:����+��9�u|\�D��08�h�A!����
D��Ĭ���<��Xl��w�/~�x��9���lx��Rn��#�^����<��ZR1��[���w�3�=���R�M��N��}m�V�IF�V��2S�¢
���#�Sz���Į�ڂ)�k���4����v�y��*����1�k�=R��M)W��$������f2d!s2��F�30�|4��H�q�4�^�W�u�tY��NGk���qR������biÚ~Q=�7 ��|��,;��d�?�HYx�L�����*��Yu�^0���nF6���u�=*G:!�T��m����+�vbHK� ���
��1K(>,����p��?�X��!U��+��Rv�Ke�"L�j�����o���#��%�>��SG7�������^�&�����î? �˕O �����:_#!�&&A��~�s���FO�;S��#XȗH!+��ۙg9>�l^�ۅux�X��S6�JmHzW���9�A֜�q��nJ�(-.f��W1���SX \qtRGFTMr R"�I�?+e�����)D��4kރG��l*����N@b\���z7�F�u{2T���SY܊��,3���<^�<�=8?ٵ�6���:'w%�׀��R�j����z�K��n�UN檱���B9�(F�/r�s�=c ���q�vp��j����$�"蒽��r���gH��`��=9��I�r��lǩ׻!��5u4�}��@W��E[ a�]����
�g,Z�<�<�#a�˄z0�w�c�f:�Y��ITd@�t�]p��c��at^.W]Vd�DUgzb�rZv�k���B����Q��	� z��4�8�Ѩ-��s�A���NI�JN�2�t��n{��4��:�$g/�/�����S���/K)�ط��ɒ�I�X�(��{�(�|*�c����N @���d���\� �`)�єW�� �m�zS�F������_r��E��	I����HZ���E+6�j�xe�X���	)�97�a>E!dH�#����O�������C�sV�!�����'�A>Fڒ�i|G3h�u�)�r��+��[��Hn(��5Tz��"[�_~�#�l��eh��Oϣ0��.��ȇ�EgG9���8b������6|����c������o!�	�ml=*�l��|��d9����*�?��B����@��6�:tK'����/��g�����j'Dݢ��l�	�iO��;I�o�Qy6�J ��ڽ���Ϛ���X�Ψo:��>��;�r5д vT.��������c>p^$!���U{�z3�f+��m�(�{��D�뱺��t��b�����:E�8�9�)��GHW��h��� yE�<A�⪙��&�Qb��dWS�Ԃ�x1*D�	��zHCa��̖�o�C�'j, ��}�A;
�G�7ub�͓�2�!�}l��!�h��{_�v!��-�T M�~�zLXʯR��o�$�W�s������;��J@1�o͜���l~�Iu���aѽ�At���S���7������E��Ѳ&�[��ꝥ4C���Ϙ~Hj�L��5R�E��'s��9��}���a3���%��|��<k<ǯ ��'��GJ�0Јf�	�;I@peTj*z1��iA-��g3el�7�o'�C5�1�/M������}
g=�!K����_��e])����*�aw�@�"�߷�"d���u��e0=�pKF��iR��F4mEw��6bG�_�<�Eӏ�98uGj����瓲�|�G�?N^�Dz��Ʈ�X���;�!0�(&i��p��$V�'+�+&�$��?w�]�_�q�X�Y�ϔx��T�|;����97�j��{
 [\��K�}�D�\^�·s;��U+�j�W(ȥ[�c`�� �9�{����o�?6��m9��;�EE�1H:��/:�e��$���`�=y�[�qs)Eи>�����vX�TK�x�y��Lꚕ$ތ�X(<�i`ti����6���ļ�2v��q��gaq�~���߹�O�/E�w(��x�6����q1y���{9�AѤL�1����~�Nm�i�0n빊�����!O�Q���l�C�R�5;�|��#�g��*�b ��Ӧ <ȋ�+�cj:��C�k��~��9U��ql?�k�A!	�|9�����3B S�{g<�B3ҷ�Z��
�]6`k���ߛ7�7��^������}��&+�r�1I2!@�a8�,��彔��%
!&�U'"g������2�O��bok��:d��$g�l�5��Փu��l܀�����,G�XEcuĮy�97T,� ����	�K~��/�U����}&`M�Lw8o�Q����q�k�C���fh�b8߈h�/}~fQ����Ch���qMdڏ���i���g{�>s��[+��&���~��m���'�w�3;2� �O���|x�[��$��qI�B/��M�.�o��	i��+�
�=�w��mXƴ}T��4�4"m8 �s�v�e�䋓�C��}2D�1q[$�4<e:|G���4�'��G���0��s���҉����*��l�`�ἵ�����,�/*P@&���=��7h�"���[�0����چON��εע"���6��3kO��s�)K�:Az%uw�>4PsY� -�4��gS�R嚇h�G����P%$b�tG!�d��Q<5�qϵ�����}�N�pΏ��R��+��s���le�+����J�cg��2x��#�9Vw�Q�P�%(P���|3��ZL��V� p�zegQ�������:/&N�P�@�����k��9�5���[M�ґ�z�画"��������� \����y�����(`y�kw����=���4 ?�Aq��^��N��(�g�$~O !.A��|�ȫ��?}��(
�'���$
yP�AG��� _�Wʗ�sB��Ȅ�s�A���ZY/���th\t��p��.�RU�,��~&�@۝>�QޯB���+_��j�􋶶,�� �_ͭ�x M�x���P��8������c�Wg�J���c��]q�q0�Z�@�o�mA�!\�7�w�2D�Ef������1x�\8v�S6]��_�1롲ӂN����+�nq�]7�G?]y�ea�2��F�i�V��������Q�;�A#F̢�X�l~�-���f+�p��y��`8����,����Jd9rڡ]�3�U���������˫�`�%@�4@���+a����+��l��QT@BB�Tbң��nQ��	(�0���t���@:%�������	��?�5~>>���y������\׹�6L��ܚ�F�{������F�;�E.�Ҥ�2����Aӵ)c7	K�_�ޝ�ނv�/B���.����C2�o e�N�OE-��<����|r+i��d�t$���h+]�
Tޘ�LS5�e�	�#�����":ͼ���u�p�c��Ai���U��u� ����:�8����I�U!�&��<��2><��=��ΞR�T���)�����O�\b���t"����RƟ����f�0}�~}��Y�O��bl�(5�_�^A��׀NB(^�n7��IO��xV�!����Zb�����H�Z(�~W�[���S���X��4���#���g�ZC����:c��Z_j�v����#VOfҚ�Wu+�i��Z�y���BkZ
4c;/@�5���M�l��dM_?�����Z�Oڞ�ƝD����a�%'�����Y�<w5~sxp�rQ;2�]b��ԕ��(&���������Z ��ꦜ�=i�%��H"��)�@�6�<�Y��cܹ�YJ��a2N+	�@hje��	��5����|Q�v���Ծ��\�3��6�������F������� �b^�N�}�c��r�%(T�F�S�2?���p�d(�U�����&,��]%�TM��1r�H�*��Y�����S��?Ͽ�0x'2"5"Tv�l.uN���3��2�l�S	/�4�j��$B52+��ƫ�WP--�*�<lM:��TJ��F�>��۴���<������G�?Rc03���Dx-�ڑT�,@2io՞�Q����|�3٠
,{<���Y `{�����V_�K��mK�)z'�����^�Ynb�\��eh.�����Ͳw��oJ�.���P�/gz�c�n������Z�[���B��O�k���D~A$�"���ߴ6�T�V�������1��bxɅ�g�_���	9�qў ���V��aܭ$�m�P�Jz��CZ�e�?�|վG�9@����ڿ�)���Y�{�U{�s\e�X)��_l��g����l6�?d�}(�r�u��C��nI�D�@�gB!��$��^ą��)�u9�Λ�U�n�q�8��9���}�2�����������V�N�����g��=rmJO����~6�}h�<�0��ՠI��a���鏾�We~�o �b���s�grǕd��v�j+h8�;�M��K ��.���4r��\a}��������h��0������wcJ�﨩�1��ZP+
 ��07�8�Y 5��*�ӕ?�c�B�g��qغy���g��C�b�G�w{��ŋ�(N�� >�����xky��&�)!?�7/���u���xK��*m�q��;�xRN����b9�& �؀p��Qy��gd���-�pU3�o2�Dwq#��A�4h�*xͰK�j�K�H8eUl�c�������/�ٯ^�I����ڨ+��qg�Riy��d�:�*�S&{�4T��%i���dc�V����Yܾ����t�����.��_ĭ� �]�������Sܷ�⡕��`�r����3�7��sF��G�ī�]N�r�.�8L���96��P�>Q˘�w�F��S�)���'�G�X;�ȝ�̛>�c}�A� �Wod0�2$���tՊǨ����P��ٖ*�Z�WP�#
�d^b�2�X���ywQgw��9����b�|]�Y�G'��O�Ҹd��`9wy���AhH���z���-��#O%��j�Q�	��wd�恝��=3P?���ߟz��~�i��˓��7�j�.��tz����`��SБ���RQ(�����8uԗJG�k�V��(���k�GHk�B�R��A�S�K�/�:�+b��	��$ݨ�|u�ʀ#@��<����/�	$]<MQ��W��(����9���y��Z���.�,ظ�j��4E�з�U�d������,'K�d�@3ɲJ��r;yB�mPYͯ�����r�Ak� L�@���� �y��҅zqQ�gY'�W�U=3�s��'/:d�d ���H�}����Qg��:�=g�'I-(EC��
�'�o'�X�rVg�Z�z/�ܩ�1n�@"��7a8J�C�0?���c�nfx��� jƭ�Ϻ�뼨�N|�Y�<��5[���zJ��e#����ΰ�U�ԋC��l��Mx��a���+�;T�4���%�"��OJ0�zi5I]�8�-<���Qm�+�~�*�y�9��tjGFJ���V�TT�Ε z�t�ڶ��%([;����͐Ӥe*�������¾��x�l��]:_d3�h��nJ���=qt�|ч�v�	pV����~���8���K�7Pˡ�(�H�r�Dsz7[o�o����9������7�o���{Û����J��i�%p����~,i-�Y�V�Zgo��X���i;�4Ǌ"\�]��o
-zV�v�U�P��Ky��ר1(S\����w�#/�m���sBM���F&\F�7/n�z�q
���?1�K�"]x0�]'���:ێ�18
t��i�݀�Q��֤�f|�d�ρ�y�z�����pϬ�p�rY#�
��� =h+�r�?��>e�A�Eb�_+���[!X����(�Q�|t{c�M���W�s��ީr�5�47a[��7�YW��%P��\ϒ������gu;��ʬI=��[����B�uB�C(�W��o�S�>�X�Jvf����7�7���`#���)�ה-�r|0��T��3�+���~�ʕv�0�g�?j�:�D�/?�{:,^4?Z�b��r�
j����+�w�]s]D�=$���.��,Ω�x���l�([r��W���eof�p�� �,m4@���Ҝ}��r�c��yc��|��Ů��k��Q�����F��s�_������ͣz��h��L�`�'}�_������w�P�B'�JK�vs
~N���7��6P�~��Lն�r�ؠ����3ǡ�>cPh�t��>���FN@��@ϯ�W19*عe�~�B�溝�����>���;n�W���B��":�;u�[��4z
d�ק\��t����E^}�pT���-˗d��ه�o/��1�����ڗ�jj��,���l"�VpV�{f+�@K����S�Lx{�F���!��?[_����AEBrz36~|���_��,U-�60�G|Z{�&�����Hu������4J�U
<w)nt���wE��6��v��)�i:�L98�4H�"�E��[U��}&)�u����#:�J6\�I7g�^�NUr�b��z�ι�����~�%*���I�����7���w:�)9���e:	���a��Z�s|`+�1�&#C���r�1��vMr&;�F�u�����H�����c�Ab|F37]���u�ˇ�,`c�Y�Ot��]<{��g�Md��8�MRN��i��6�b}���s ��`9�˞��ǜswu��Fmh�q��7+Vڢ%5�]����t���,�9�x@y�>D�44r@��P�<&���b\�3���p��S]�'�C��Zj�|�
�BC���Pt��*��o޼G��2�����{4���@������@���=d�{�B]����� G_�G~�w��6ڋu�8h/�!�5�9G��J�-�H�E���͆~A'�$_���w��ܢ���YC���s�T�.�B'T��Fc�T/hN�����6��dqS,M�=J��Rs�}�S�C���oC6� A����kt����q�4k	ȳ���/�A�N�#.�y!�!*Z��e��oŠ��*)��j�����U�L���
���,G����j��_���9���c�M_N?�l���5������慞�
[�����x+�ø q�H�J�+�]�C�[�?�>�S$�x8&;��9 �{�O~�k��st�����C��U;�X[�irV�a	�&�:)IŚ�',�ӝ) �`�`����7�~������f�Z�.'�*��-̮�%��^2���D�I��	��'J>�{U@[�#[tY{�YWɌ��cc���3�܍_���U�77�v9�����C�F̯��?ň�H�D�ؓ����6�����2�X�7�Glj�$=�J��c������&Oy���Δ��v:i����ؖ 涭�7^\|�c�Tc����hY���N�y�ޚ���!��{�0�Č��T85k�S������4�[S����W��2�qe���;g2MsV�!g���D1��/��X�ݞfpK����B��@���u�pv5R�$��	oC�����~�;NT�_v�_LG�[�]�ڄy�n%��r�e�Z���8J|�֬�a0��>q!�h�A��@lu5����|�+d;��^�j��K�:�?嚎�8ϊ��4��\�s]D%�@��[�O�^c�ѓ�Jn<���ǎ�Ue-�h�XKX�d�;��]V��nQA���݋Po{�#d�IQ��\�HӐ����N��x�;��{V��G'�l�_M�}�8dQ7��V��(�#��:�
��y�z� �Ce�:I�L�����7��9H��[-�L�J^D�s���E4���ȄTm��9�6�Ր_���qg���j|�Z�f�9�Ǟ<N�Ͻr�6��o��&�7���h��G@4��@�&�72^��L�����>�[|Ũ���u��#A�Bm�C'���s��P���Rx������WRKTT��AH��\�7�wD��|������[��q�k	=���tb볭PSU|pj����Aє�DNѭ��l���-��b©����i(2�d�䛓d4�rz��\/�$ٙ�]��б˥��Լyس�C�_�-V�w���ө�����_\�o������Z�)M7J��*�±.1ޑ�sV ���B�rk^b�k�u�а��3On< 
:�	Vv-� �M�pFyn��J��z��4��)���t�K��vVu7�؉��	6@=�$�ѡ����]�q�BӾ�"�����N�=-L���K�73�^	�I�?��YE��h?�*^���'�WlNM\P�v e
��xV��� xA��l���L�L�9rV��WR8�9��ٜx��(�p ���7y�5l�X;�Tz�Y`�'�#�iM�d�{�.Ʀ\���[��^�A�Jܑ�	ky�h��Ui'*,�Gp�GlÜ�^1 �
)N�c�m4�;m-����˥BXήM�*��I�Rc�4
����IO�� �ܙ��Ìu�b�ⵠ�i���ZǊW2(V���s�oO(�#🣁�����5�)j���J����h.q����NA�qy��au���r��҄��"u��еJ�8��Ϻ/H�>h���\m ��V��M�u��?�R��5W{��Amꢊ �m�����ѡ"���&���[(���4��z�W�jD�S'ߙ0��?���#ѧ�*�����3��4���-���N��C��(>�k�IQ� Rq�h�_$�T�_�����;|~LS"�J�Ԭ2���N���Pa��o��(grϡւ���ҌM@������Vl�u=�ϵ+�+�;�sbW�^k\<}j��p��$Yi��Ý���f@!�)1ϟx�U%��K5M�:O
5����{Q�Я
0Ϥ8� ������K��q�z�.��z�	�o��U�^����Α��QG�r�S��xw��Q�򑴉�jH��F���4�8����{�5Y���C�H�ȼ�����r�1�u�x;�Ԕ�p��@L�5g����fEN �-�9�x�Eޭו�	
A�� ��wX��5���IW��><=�_�@~DyodC߬Hj_}ؖE\��r3 ~5
�{ȏ���K.��,�e[[gsm�܉�:W�T�{y�i��΀hM��H{0;`N�z�?�=A��ʗm��=՛�˼��7�Y4���;� ��t]� ��P��l�|.f	� C�"a�p��q�3U�����ܸ�*}�䓸!ֆ�۲��u�2�W�	W>U�X,�f8U�m�����Q8�u2�4�	�>�sh#�u��"��f�V`#_��}Y'b�B����ͥKO>	�4/x�F���i�������1˥��]oD�mڿ�R}�B#J�A;0��I�2h8	o�u��ݕ{�����>r���C2�=U� m y�5����la����"�/����l�tO�����c��F�O���d���=Y�U�^���d���ś���L�[�h���h�������^�|D�s`��_�3����S�^�#Ƶ�
������1��}j�;� ��_�g�z�n�1�&�4g�k���y�b�~�[^@M>�o�hX+G�K��L��	Ch�:�v�P}�#�G���n�r$�EQ�zW�9���f���e�껝�kT�������
�������f�c��i��4r/RX�i����w��?�^�J���"ŉ�P�s�M]���,5"�vrE��Q�gE��)���T�;Ͷ%�i��bsr3ǐ(���X�����M��Xe�!�x�R|��i%\J��M���6�k�M��ƌhב�p��W)O7�nU��j�!��w�Xz�Ƥ�����{DÇ��s�M��n{�-���έ��ͥ4�m����4�.��r!	�³0�⫔�Y\��\�zkrp);�m�i�'a��x,Q�v�ʛ�6���3N�(�EZ��2��嗮��Z�L}o�����|���fG�����k���^N?�~������i{@H,j�^ѐ�\�� {��	ل�.���5~������6��| �se����N�"E��]��7?��R75���KYTﳥ�dT{���<�^�|t�ޣ�����}E��>�.3霠�ND���.��ud���ӊ[��
S�o���&�����J���A�iz�q���.�Yb��E3���U��x�q�5v���n͠o��"vפ�g�l��L����3x|�L���=�����>��j���M�Ox�j�|��[,���0ˇ�@��������գ�kY���n��"��+�Ir�`��f-M��6��[4�[�b��p�N=�h�c,������^1[U�/�౲lSC�nxu:���Δ��%�Hd���k~S_+56FO�{;�.
x���j�Zڵ����[|�MŌ�G�A�ԙA��T��h�j{9�ٲ�sW�ј��#5�����˓Ak��FH7!d����Sf��ؒĴw�Pii�״��R��^H��bS{��2��N��^a̬۵��ISR|6q{'f��>3��5Z~�E��gĲ;��'!AX�Q�.g�"�Cѽ�y_o�2A�]z�Y��ê:=)Ƿ��HZ)\t.��]w�j��Ux�lA��6��ڢv���`����{˫��N��E�"5�r�j��ΡKT�C�$�n�����XJf���)x��A�!���e�y�o�l�E�^5a��6~	����,1{�L\�̗�0�^��ܳ�s��&?'c�k/)_��5Y)"/�Sc�澛�k)_��nw��)�e���eB�|���߰�Ö[�7"cq0e���6^��(p	�5֌D*�U���ټ/�Y�&&��S�Ӿ������+��;Yhqk��J��U<��}�	�
ꎘ�͢j��`41��PG�\2�l}��ꑧ��bVRR%8[IHˊ��P��-��t�O]�7�X�(wB��	X��(�|;��L8��jDj}{��_��QҎc�f;'��6%����X0}����H�{T�����]IERm��q�Y!Z��\L�ދ�tk��7����k1CΫ})��t-�])��D�9���Mق$�ʹ2;�׌V$$��On�B��*�I�����̺��J���Dަ%#OA��0�)���Z�_~~����K�M׬Q՘��d}2f��h�PR@zĈL��S]7� ��fH�M��PtVN�`��dt�r�AЄ���Tӗ5�	K
IX��H����Nd4j��5�H�[�+�k���`�l���������6��7��3��������S�~aB���@M|��a��C&%iH�AFw�ktp�}ME�LGK�ь����H��Z8I�_��@����d���
�&���5�Xqp�ĸt �ɘ����*�:�(ɫ�rV����$ܧ�u3�Й>А&�H�����[����Wlg@�"J�ů���Z�o�;Oz5���l��̑�:P+̀���+է�R�+�������o7,��cmW��[������Rk��qV5Vn���+ַc�J�7a~���R�fGg5��8��e�V�HŽ"O�{E�>6$H�����<ƥ�bp+<L9@�2�H��|Fΰ�~|�sg�����T�^*U_�r�G}l�b39�aZ�|}��y�c��D��~��O�,�OHUʼ����M�qo`�.=���Ijw��M�lx��P��I�5�R��hm��u�;_ҳ�C�e�Y�:�2zq�U�J�ܳ[��3�Ec5($�|��̆��;�i<>Q��e������<Ʋа� ��J#�������ݙ2I=�Y9�_8)|}�X���X��m>����a��ӡb���_�k=W:y#����Β������<+s2Dg����*^��)�,�iz��ys�rR�7��
��$7�<�$��0E�����a�B�{�93�Ӷ���.�)�~�y��@:�F�Wِ�"ʴ%���ų�VW�]z2b�e(~�0X	{b��f=�CG�Iiܗj[�?@Ö�|rk'p��Cq%�Ls�%.�ce���5�m�Q�͜]F�@{`Q�D��f!����M�H�� �Jq��8��Y�4���Vq��a�̔[(��c��B�b����,%�U1?S�Ê-��=�[^�D��c$Zv�m�l^��ق���W��w�
��i��zhwTl�Hq��VD����裵bo��ߚ�������A�9$�&��xe�Iӛe	�,$ǵ���v��J3�|�Yi�d�aY����QR�������'��g<�p�`u�[<�2��x��n*�L�������>R+V�#�^���IF�맖/���WEC���h���%F��6C7�=U�x�F�k��r���V_����"%Ic�}K%���M,����0��g�����h�xRʟp�D~������,h��X}367���=�U>��l�����La{C��%��$�� k�ڞ~kյ��H���̋���Û$jE�}2Mǥ���K�yVIB�3KH�w����2	���^���4-��)�H���𗓫�͵^�t �>��cHL�;����D��六�@%��n�r xU��N��U����H�j���馓	��0�\t�������y��- <�K��dZ�n�A&��B�SEO3!
�K��f��˹1��GTQ�^͠Kv���?XYSCìf�'x�)rHd��\MF�;YZ'2�)��$�IZWE#���
ʯ������ڱ�A@��T���UAko�&���&0�T�OJ'���%�|�@���D���Z2�������ncO��@���u,�>������430���f�<� ["�f퍂�>��2%�R��&z���f���1+�8*�b1��e�&x��o�(����ѵ�� 9 ��r�V<�N����b�PNz�1/�l��F�O���")G��5�V	1�ra�����-��66�����Q���f�e�ϦilK�Lb��gN�����`�o���i�%��(tX5~-*�Nh؜祔;jFGo�s�GL�VOZ���0����M��pD�^Oo�M)QP#u2�B�d���=���G��M�Y�ZN~T3���<c+�:�����2j���u��5u��ݢ��$M��9���,���V���/�s��ʼx��d��,'M|��?a��e��qˬ��#��+1Ξ��$�O%Nl:�3�bȰ��)���L��Z������o�+bC�k�!e��{�C�2[�u���K��������dj}� `�גR&��@P���_=�����D�f8Ƴ�I��?] ^�;ݹM#�^�_NM��z�}�h����u>��]�� ���;CK�ήy	nzU��KKɹ�T���lx@o"l������8c��j���)@5]�7w��*lPj2���A�[�%$H��wcpԍ��D�*gŊHQ�EC�2�4��4�y�K���Z�mʣV}��q�gv�h�:)���n&�_pC�v;�,I���������D�~��/���!sXơ ��ZT��zW��'��Q��opLy�M�$��ڪ�mɧ&��g������9�3�:3լ�A�:Z�Ɏ�A����IS��
�������?P�#c�X�P�����*F)��3�Q⠌A�t����\��'�Oz�E�~����#s��N��/[i��.�mb������a��I ���@��8��hA�64�X��R�w�?'��6�u��>-����"�"R���!)uV_?;�XU��hyc� ����; )	r�j��z�X�U|���
0���#g)q�:��Qu᠂��ds�s�t�K�}b6��������|>�ݨ��a��#&�ݻ�|�u��݌����{:C�GXz"935��{0Qg@d��LYq��� �[��C�j\�)����y{����8tOǲ���*�-��<
�/Ņ���
Okm�s�f�~s�I{f��$*ͳD����o�X�[{O��k�Z�I�qE&e+(� ���xek��ޮ��N�fjG��)C�\��{�L�a�c����W�P�f������ټ��Ya�?����I��T��F+�%�'��o�]��wI��� �K�F7nO3�g��j<�z~�g�|u	�$��jR�n@{��􅅳uIne�t4u鎞+M�7�1��H�JJ��ЂD6�������;Šr��sSQ+]��E��zzڧy Ӂ�!�K=�l{�4����(����0�_�m�:����{�̈́l���v��6b4u�Ƒ�ɳIF�ע�SȊA;6s����&ᡢW�fh�3�eR��m��	w>^�DM<o�7��X=�5H����� �##[5�Z_��-<`6��΃�b��{yܔ����O�Ã��45s��*��+�*�W	j%�x����A�_DV���I�
}z�FI9��xR(��Py�um}OJ<����ܝ�	V��ßI$3��P/{��k6��҂���Z�V�N}9���vk���RD�E{�ӝ�ˠơ�
8��յ�m,��s���c�5)H!����3������w�?�E��Z[����cй�K�*��Ⱥu����)՗@�;|���9@;N��O\M
S��`Z81�ѿ���ne�����yH���_^����ޝ�����'��oSb��F��߅c�xtu�H���� ���<Q���2�5�q/y��GpD�?�}CGXÁ\�f�/.]�T����/}�#ױD�p#l�|~�^��?��w���!�,�!'ũhq�jz�]?�MR	$n�l��"(��ŀD�;��E��!�;����M@r��qѺ��&!	����ݹb!�KS_��R1�zEW͓�6�����x��������Ҿ���O�J]�rݡ@`(����bp�M�m����5�W�:�1����,�ï�>+Ǎ}D<Wd�Qj�%�n6���Q	)>ϟH�t��I��5�V�@,F�Y���d�}W�<B��a����Z����7�/�/Eh���X�)���e]�M����U d��`��SB!��s���p��<�Α��15�c�#
}R%���n��%�Q�K�e6�c��<������ ����F��&�� ���[�^P���P	8���$n��WnA:e�4eBP��c�g��S��:\������I�Yw��%�3�)��zn�q�:��K�F?3i�ё�p_����@����Ҁd�jDO��m��*B�J�w]�H�
�u���lJ�%�9G/�}��R|�H�6j�Q����.@��'����3P]w���Bͤ����M�m����	H�������x�k:��Y=���a���ݮկ��&m	I���$��������� ;�uB�E�g�3n���"�x�8�&�ۊ͝��̽
�I/��76��&D=�	L`h���nx�/#ò��x�Yp��RX��x^��oy!a���� _�����ï�a$�1��e��E]�������ޡkYx�r8�L䂵�ϼ���"�=�fҢ��L% ����ǥ��}h4�kd
}�
p����*�1ȹ�ۼ���N��禤�w�}q�Bȣ͵h.�C�fb3�����-���m��{�L ����s_�)���X��ˤ�(,n{�'!F���s�?�*�< 2�����s�@��rB�a����)������r;�u��1�W���AI`�<�XqnE4cz��t+
��M��(ΐ���"�:���!Ӆ�w�l{M����G=�м��zͣ/�Z��`����!;���f�\�����۷/�$c��E[F�Zͬ��ｕ���X���\M���X��0�!z_�<,�G��
���Q�ն���[��u����q~ SE+-����)��vG�8�ew@7G���(M�y����	?��G�V��D��f`
շL<�R9ô�yt��[���X�BE����B�����p߳�*J�8MO�{� ���b?���4���n~���]���E�CW_�HH��t4�ux]��46iw���_���E��ݭڱo����@m�q��A!�Ju�� �apT7�ϼD�"���e��*�4��>g�r#�l�Ƈ��D�}L�nM�;�������S�J�̿�v3��7����'����mE4���	ܸۊ�5��Y��X$Z�"^�� ����9X�;��j^C�����g,o�3�jz!�G�<���ěkj���S`��Vc��.�dR3�:=��~;/Uְ��Dߥ�Rk<�6�h�I(aчj��CH,��pm$17�{��1v��"J2���	��@���O�*DB���"3{����^)�|�����w}��QK2+]r�d ��|)���'�$Xk�F����s���]��b���/D��d'�}a��\{�s�B̉�`/�Q���E�U��v�/�f�:���2*�/�����̪�$�b��j�z� (|2������'$W�����Y�����gI]�S� 6a�A)<�`��l*�s>u!8р=������g����R� ��Z0ݶ9Ė�I�>�n_��L̑F�Xy���E	��Q���ERK�^y�����1>����x��}���\� t6�H�pY�^�o�i�����1_w�
J[Bds)�AL�k�Vp5A�([��#�1�`�a5�|	���4���K��B�n:7%5X��\�6!z�I���o��R�f�K�/�z��U�1ձ��y��kH
�F�����DO3!�~�?���B5a���$s�V�+�J�����|�K897H���`Hy����g��c�Ck�H���aFt"I�w6���K�E����hSn-��f{�̟H7����]�y��*�9}�X�[�;K��yo�����#^�f��6,)��
�Nto�բ_G�����s2��n�ܪ.e%ve"ڛdΔ�c��n�����}�h�a�R���=Хf߾�'��ǹ�T���s�{�BV��e�/����[}3H ,��5�R"^���6⿗l�ac{w��M�gOg;�����@��U�)��<Q'H][daI �"�	l) �u�HY@)�m�3B}��]�E�?wPwI�`7���9�q���@l�ʸ���{ ��4�52D�Xʰ�Jo�B����_o��"�Q`:s,%����W�\�)���>�U��Jl�u�g[�]�����9;���Ї7��P/�-z���~	'�Jਿ�+T���b#�s�p�$�" �<q�/�}�l5�j4`-���Eͯ�v��E���7:�	�.'z��k���;��h�{�p	�L����D�p�'��PwAg�D���p�H�eM�ʟ����	������3z�f1�����i�����)Hs�����}.Z�
�G R��x-ʶl��Q͂?�����~�$�̒4~dk�
0W�{*��g{S��_�tR�\��ҵ�"K��'���.�GU9�K��FǦ������+o�<�P ��<�ߏ Yo~0�H�b�¼��u t8:Aq4�!υJ�]G�"�6�Q��w ��0��2T���?ǔ�K�[E��|�,�.�A��m�R{�b[�٣֌S'����
�����f��[���Y
"�Q����`�Bw�C,�N�Ub����A��#��e�΍+Pl��_F~/�e���&�+~�e�6����	ڐ��ֻ���A�$�C��w�!X
�Ow�!Ȫ�Ofa��\(���008��4��ʠ��/�aQ]�0j���:��Y`�EU\O�����o�K��%4��jY��Ю�� �C-��W�c���篻k�܄�?5v�ߠ�_��dyyyP��Ax�t�r�J3�N�N<
�("_>�)4�1� ���r�׋^�>Pu�t�{��m$�D7��t��,�
ku���KAx6Z�J�l�e-h1�F��K�nJx��S􍵃��x�1�R�Y�Ϗ�H*���:}.(�"W)���'WT/�⽗_�+(�7��;(Ù�V�a?���1$�r ��v�)� N���S^�1i���a������
�%0u���lH�@��#9(cT@c���7/0+CI�T4���TA#����F>*������6�s P��N����
k^�n|��j�y��h�;��t!S�7v6�NF��]u[���2�|-�Kx}2v��t��+���%�.��c��rN͊g�+~�bv�L<��i�U����'�10c$�à��nd���{�`^����Fx/R���Qm���������8Uj��d}r��l�'�!4�R:87�G�� ��@~h-?d��/>�G���N�����P:�ZP&���R���ʃ�ñ���L̖��ҁ1>M��,d^|�^q�>?��饿�I����]���
:�دb���z���fI3����Zm��+��R!�<��i̹���38q�����5�`����$�F`�6�<�4`�G	���s�%�i��#���Y��+�i@�r1{р��i<`�9�C,cvZlFα���`ʍ�O��`�<��R�����1����X����Ď�������]yx��~Љ\CC3+�B���~?���l��(���-t�^$�q��26��$qj2�|����Н������U�YU����bW��S ���k� �\�G<,����@�V����]K\JXe�������lkx�ݦN��m��#��o�¶��!_��~��ߡ�6w̕�"���^�%B���KDe��B�����6bٓ�u#�n�I�����7��M�x(.QZK�V ��c�c�Rb:21�Ŵ�0�9�0�1�
�� V�t�� XH�@��隞6_W=ꡰ�!s8�&�����zu)��Y�d�����y�}����K���q0G��F�i�����˚x;QkhH(0pQ91��T�E3t�{{�Iof�Y'տ�˻
b�2��l�M <��Rx�p����ȏu5��sa��>�q{��:1@��Fpąo=j�L48N�̈́��ɰݗ�a?ʔ��;�۷I@�2�Bz�{-��, Pm��°B;�v���PK��'����2�L�ߔ7����I]��9�O�m~�MQ���
Ȕ�������5�v��(�AĮ���t���������D�}��"L�s��?�a�T�g��y���6rfm7S���8��н������@IC�Sص�&j��{^;!Ak�4.c싸Q�.5�ʥ�2����>���'��_�h�K),���hM�U���caa �B�\E355��K|=�r؇j�&챞��ץ��qV~����m,&�峠��H�wZ�ў@�Y0�'tp�å���V  ��71�m����b�}�������b��e�X��pI��6xz�3�Y�;=( ɰ��&����'u5�����|�{�L�T�lVNvPV~���n��)9��9KIb��/��8iΞ-M
X5�ǻ�	O�~@�(�Qc �fh�/���%u}���CK��'��؟���B��(i�=�YK%��Gߒ<� ���3�_qΨ$]���Ͽ��_��a<-�g,D�|��v2�f(%��FhV���L���4��&
o���v��p��OL-������k��������	WO5��G���
��;@�!d�}�0���+��7w�G��nL���) ��}����H~Ĭ�}&�m� +�����O֙�;��|r7=�߃����[S��gҝ����g�yuH;���w��aPc��R��hGP�\P9�'ђ��p�T�?��~ik�� R5#��Y(���6)��n��1B�@._-������s��X޼��^h�k����
��έ�Hl�?�p�š�6�q���-�,�����
��|O~�����U��RQ+�������>�O�`���03sU��v��;%�&
謬���1$���f*%g�l��I�2���l�Q��/��T���JI�E,�i km)HY�H{l�Q��f1�G�}�:�̦���W��W��p�W���Z-]61��-�˺r>6��	]��3�:~��ژ��ɺ�|�@����%.E��e.cj�8f�򓚞��Z���������w�E��S��x�w�ɮa�p�Ѷ��)b�l^�P�㻔��N�,h~o{��~{��u�c��ߢ-��A�Qy{��4�KS�*&���Z��*�罺��|�ث$-6�����]����V�	�D&m�Ϫ%�5��;���٘��3��RD�d{���{`�����m̐ �e[З��;�UK _��S�-�D�?e��`���U{׻-�;��;��_�5-�^Z��@��#�gۆ��z��9���qO E��q31���:1�(}�{1pPV�Q~����k���s��5�34�"��͙�7����晘K�2��	�U�	P�H�+�-�\��U"څ4�`��]0����?Vգ;�:�]y���;�+e�۫E��K���zOo7�{�f6b>>6�RZ6N{?�6mm��D�KA$����_��m�VK8�B���S�1��91�SQz��8�Y�0�h�/�A����ػK9�El��-!��1JC-D�������^�������'��	�k��	��Xz,��]�vQ���N����Xk|b+�8H%.I�١���!�;�mn��5�{�ڢe'�弊������WmL���X��-b�1��z�q��Ͳ4�Bݜ�Tk�t�{���"�%Ď�+����`�p(��N�+/=y����
�K"sx�Z��gamAs+=ͬP�R,?e%
��85��uS�d� �����	mHC�;z2�If�/>��T��52O�� ^q�R���Dȣ'h�W+�B&f3��$�.Bpj0ÉU�:�����Ɠ�x/���IV)���c5#Ҏ��,��L�p�=�!v$�;���EÚ+9�����Y��Sb��%�4C�/&d�I$Iݖ>�-͌�<~�$.��ٺ�o��$RRu^挮a�N���V�&����v��YR����[���X{��gN=p���#�o��{t�;W���1��/~v6��%��KY�IE=���SE����YR|��Ŷ%�߯�a���x�׻��oU౶dE��	e�o\YA�8a�-�N
�m��%�6���l�������A0�d��kZ�Gop�ת��c�;_no��Bn�ޞ(��r��iG�oEN��]�X�����{F5��{�l�� @QA���Ԁ
� R�lPP@z%�"JUz
Ҥ��ҤF���%��I�L֊���/w�q�9�u���aε��~O�%3�V:��^�+��W� �E�;z�2�����^)��E�($U6�d�p�<?��[�����z:��B�i�8�i�ɰ�#��Ļ;V�$0�RÃ1�&G��c|��y٫CD61�����>�W��x�x���U�9��~ʨe��@Z��{�[w0�S�uhŏ��-Ĕ����W����&�N���4�wZN�5�ٹL��IWz-x��˝����:R9ݭ���Y9�[�s�qx)� pnÆ����1eh�l����Y��;7�1�MLD�����iEW^���)6xx/�Ǫ�� ��1f��$_k:,5c�J3�X`��dC���uA0~�f��'���5˔�^�(�
~}�T�wbt�����*}�o�(��>&~�\�6m��O�F��|,�I$��]�5�6��sq�Գ	���AdO�ȞH\�Df�L���TmR��gu����9�^���j�H��V&Z*�Z9E���5KT�o���v���s÷'��F���rЦ�~��Km��#���؄�	g�]�r�bz�3��ݢ!\M[s�$��x�ڸ����ƪT�#N<)���&��Z<o�Oc�Ή��x���,��!���Sո���gS�۵����F���'���i��e��H��=�]zm�[�".PQ��u�j�m喴w=GrB�taNu����R�s�p^BGG����Š����D� lv�5r6ۮe7+�}?�\��U� .���:F��c�=�:$�V���\���9gүHݻ�ԡp]ʠ����^�-�������������<N�Qj�3{�āv0j%���Lw8��,E����k#��<�ڌO-t��d;M�g�������\�}hU��PI��M-}�-�D���CTBTR��wۧ^����@���]�˻3p�jRq�O���7�C,���YX9�;��h����J��a���ށz�첦;y�ȓȍAt�{G�oM	Yi�#}�'0�܉ͱ�Xn�J_�-m���k��ɗ���ʯ��{���������́�����] ��x�uQ�z�^��i�IZ���R��5��^���O�r�o^��n�(!!.n��bRb�r�N\+i)\�!��Poq/�����+��v�<.����x6�9%}M���ɊFΤ������L|��\�U����|yNηF�ފN:���Mߛ^M�V��KZ�Ul����i��R⮽������/К�e���(���c��F@����a����,b�M��O��_�
Z)c)�h��ώ4�1����',�Z�C����~m��<y^}�A[��g�bjgP<�k/��Gu���9'�#eVti�q*�0���Tz��娑��(qq�,�j��%Wp��ZKx1^6��LA��c�l��8��G�%�M��%k��,Eg���ģw����Q�P�?�N$(́RoƆ��H_�|������:�w�@�ǽ�?�׈KU`�}��|1�T�)��k�' �k[�Ln<k����$�3�q� �hPE�%σ���)��.��Ew�p?C��*�"3�b� ���I
��oo��?F����R���KdߓA�3*�����(�/{q�X|��2����[���Nb���F�㼧�:̶5;t�%*�Rc4�H˗��SQs� �i�8� � ���K�5E����e4x�����`Ve�L�x����󹛔��·ʰ*xL; �',����)m:���|���	��S:�$�����9\���|���M3�J`띯��]��!U�L�qc�9^i����d�[�T_)\�x_�(��41�<�{�R|�޺�b�Yg�����)3S1�����F2�%�����c!IV͇'2�=1��(���ܚ�.t�܋�~�WDq�៧6�聘�&���)�5b�5�+��>��	g��D*^����N_̜���-?6z�Tj�6��K��6zl�W���Cm�m�ASW�
�a����R�����8�#w�e��+�p�i��
�aH�!�\�M��E�����2^b�q=��jyw��d�F5.��ᖢ�	0���|�IM.� ��ݞ��qS� ��'_eu���i�PQӾ�E���x��h;k�@��}�p�G�oIa��/]C�i)r�$�w���a_a�o��Oj�7�;�C����x)�����=��|�p80���n�ϡa��y��Å��ӹ�Ug-���1��Hi�U�xq�#bGqr��4�\&I�`���:��Y<��	�@�x�1SPx��?ݝVp���OR��/%�ꇿ=��Y���p1�����w��[_�A�U��V��jwZ�h��a%��FI��i�?K�&@����0��c��Z=�Q���1F-_�kP�Q��3�9g�y�F�qj��k:(~�Sʆ��e׾f�p����v�=ONL�PLy�
�#�;��܉3�8�K�&��:�o�<E�~��@�>V/�3<tB̶>������V��@�D�X$%�=gH�'1�wW�ҫ�����7&�Q�nJ;"1�u<����o/�3��*
87���T� AV>I��&�n�vf ��Zs��&�s�GTxZƽov�;b|@�D��"A���V�ݗ�.��Il]��?H*eg�� ��$ۃԪͭ� ��b����"��{/9c���[J�&d� �k��c�ŢV��"i���s����q�
ց3y�u�WW�b���]2"^J*�}�B��x |A*���j
P3׵����U�=W��/&�PD^` ��1�Qr�c�`��e�R~6�׃.������<�:��N� ��0�X��$��=����E�`����-RMF�>��e��e�;���>���o��7�x������D��= jG3O���Xލ�,nM�C�;�ңOCF�����q�A����#��:W��fE�J� �n�޿(޹�Fo8*>1�e�tĔ�z���ѥi�^kq0O���9�,��׮VώЃV~�(;����o���$����>��R�^INO�`��	�re���b�!�7G%�X�Nk��c#����.K[����{(��I�)T�H�	|�W���G�5s�n���kWD�C�Q��l��%¢��6��D=����,1ϓ��Lb�\����.m��'�����b����z�����q���B��{^+�L!�f�[;a53Fb�w������-����'x�X
����Y�1-����	����#����ǚ�&Q��ή�[c�^f�}�=�Dt�������z����>�w\�@�l��ʭ��хݿ�u�I�h=���=X�6��!(�
�'"κ�����Ou�f4�me�xj�jrNxX�$	�g�d	J�Mލd�z&8>Nc9���m����*�A={���W~��4Һ��[�ϔޖ���
E�.����'r���D�+9?4�'x�>"4^�z�+���ՌJ���*7��,f�������~D��^ޔ9q�&�%0�6%qk����b�]��?�;Fװ:ZVcR ����ό�QI�E0r4����Kĥ̲q���Ʀ���f��@�
%N1��Xj0�AXS�����Q��˸�;�{"7J����e�[ص�C芣6(Á �ZM$�z?�A�8֧6�:�
�B����ȯ�UU[�C��<�l��R� �F���)��e��H�������l���ǚ*$rt
��l���.)_?gO�~j������?����4�Fh}]R�#:r�,�d�|,H,}0���K���Á )H` �i{�LD���VT2�B��Y�Z�9H��5)�왉C0���7�  �?�@�/����3o�����U���6�3q�s]bI~Q�t�N�כ ��9'$|���+�����=���i�e�:7ڸ+g	�|�}��D���$/x�_�*x���鍻���K�WYq����F�~1�j��`&�G@�y� g���B�	$y��w�4�3�޼|�zF��F~�YP��"�Ӷ�9����^�8������G,V�ђ=�xe�8��J�ʘ��E~��e�-]M��$�'s����x��U����	�����h�	I�y���<g��#���H?��i�]��Dfr��ߏ�|HX��c�99���TrȣU���I�s/n�y|a�t�� ��+E�i̘mL��4#��$D�Q�.+�3��xQ�yD�s�ŽpM%���#�j�~d7He�
����L���˕�bE�/��A�xs�dt����_��8�����u�j�
�A1��6�Kժ~\
�Ge_P���П�I�u�ӗ��d���-ε�BC[�������32q������Ik�5�棟�_��*=�2M������z�{^W�
�L8B�l��[�ohNc��8q?��P���'ήD��Ł��K�I�]�{7��<�2�#v�ǡ��W�^�{A��!b�Ž��:��)q�d�����}�v w��������vH^����~�G��š+{c�h�x隐�f��X�цT:������Z��\t�$ x!���qt�̪�E&�����>�ٽX|����|lkU�0zV���^�Qk������T�*��ڶ�b�~��.����:�=߭m.������T����ߍ�۶�"�Uw���UO#Ok3�����r�Zک�n��|�r$�{g۸��.l9g,�M�A�����og��9 �m�X���jх�ΥY�o�v	�;���g�u8�-z�'�miH�ZXt�u�bd��﷋��+��Л�d!��~��&�%3�0ӹ�&�)��NJ�z�-�V�� �������&y�9�T�`�p{��e�����}(����Ƨ=c�^a��x}*�,��췿:��͂�`�q�Cۙu7�g:1�6:��*%R�߮��T�F'5k��ƭǶ#ˬ��G\T�A�|7�]9���'t|���=�V�����\x��f���h����w�-��jpe��y�oj ���0�"�H�p����OvϽ��|0��/ �$z�D� 7��+���(cM�����ڌ��	��[_���vmO!$�y3�8 �s��&�k�w|��Oj��V9!]��^���^ 
�wiL+�����O�)oW�M�]Ew�\��l�H�
�۰��^��73�+�_xw��e�v��GЬ�>�ˋ���|������4U/�	�v�4���q�v���QoM��"՜j�v����Ey9�@2�`b�N�6�/�Wؕ0��ۅp����e�0+)z��m��R�So�Y1߅�ϓ(�H����b-C$ìQ�����W*�^2��\�|؋�};;ۈӺ������og�ϬE��v"|�����s4(za1B��_ۼ㝁(X�mM0Ӷr�����z�PN������}�]��ʳ��Ib��(($�l�g���S�f��w(��N3�d���|e��$ݶ�v|��a�1V�
e��v\�H��kdq�F�>���7�%�O3𩹒6�9����6����� j�H� ��\�]19+�3�=1��Q`D����<��)��G΍}^���Z�ˌWvJ��<l�|�������R�S@����ԕ�F�h	]V�O9���I��_&L
n�)��o#�Z9C�۞(�o���:�t�����?����X8�C\�B���*ǧ	M~Iq0��s(m�[��	$gr���D#��u��'��B-v=��A����$m,
�E��֝�h�������O��?���:Õh@͔��'%Ň�d����.��p��u!ď��m��V���J%�;��|E��HZ+��al�������KC{2�"��Ti�����(�B���龾d�G�k槴��]��ׄB��}��q<{­!���ֽ{��[�zA����-ZE��V�#6
�N2��:z��Ղ��N�W.�a�X�T�Zd�ހ�\{2o�� L���E
�S���I�8�w�Wˁm�+����ś��GS��H�!����H�O�ev{�RӠ���|%����6s��m�!�ߕd��Z��6ז�]�;B��������5�5Z]Vf�:�*����8-Jf�7%�!R�=�2*��p���Gޅ�
��|�K�8�MR�ո%��b{6���4|�X����T�3v�'�|� �W�u>�ֶ��t��t��÷C1��glc�_[������ٕ��_�W�Ƹ�Nc��H�\��5�xWB�����j�-��~i왡��V���@C�BX!��?O��ۋU�n�k=��3�����Q�wJcr�����~�0��^����C����и�����Ɓ�4�am�<,����s�]_O�b_?]Rrr�e�͙�`5�Y�U+O��W6�����F�Wa�6)>>���	��z��}���O䫨$J���=��>��ĝ�F� E�E��{j������m��5$�țPL1��<�i�;h�;s.�;�$*C�ĝy%� �[���]Ʋ��b�i��G���B��\7�"p=�����C,SUЗ�?��	�Q�A=�?I�W\�
kޜB�v>�լZ��)���\�1��h�D%o��,��L^Z��/:5F@���8e�钬���d�mtŪW�A_�� Dmz��%�H��\$~G��+C?�y����_�Pd?�[E��[�[��%|��c�QG�&�謌<�P\�j��5�&.W���"�zƥ(�Tl�zpf�,y|�#��v��|=RG %��9.D��a�6�=M�{f��:ч��t��Y���z�o��ѭ'�O���L��S\ց���%�]������R���'?�F?2�i�����W�x���B��w`�!���yp��c2��3d�\�|e��A�������j�'Ő.��a�����g�uBg�(.y�s�H��B���rH�=66i��`i�&[MX$��)��4<��"@E��Sh�����b�R0�\An�
�9�u��WI�m1������{)*Vԩ3MiR~���o��H���1�hx�p��O�,ؚ��V���a]�����!�\t��v�W���q��K�T�w)(h�y��ٌ��P#̮��Qj*��̀�j���RH��0���[�_���a�?���f�r�*�G�e&��VIr>�~�6$�F����� ���L�E
�G2�4���x�w����h�����Ϟ1��I5�̻ce����h?5Q���B#M��E�ꣳ�>]�eF�P����E����~���1�����'!.<�&HD�«3-0�?	�X���{�&7&lt��5�O��5���]o	2��N>���&�_7Q�d��>����`� 1J<O��9�(S�ɤ�$�>yÀ�!��gv�h:��"�յ��=Êu6�����Ո�N2������N�Q�nT%}����<����q�>q8(�ʐG�l	ce����&7��Jn�΀��e!S��ۂ���W�2�INe�^� �t_�K�2`�_v�yE3�M>Ђ���H�v�0�������(x�268Є�� �螀�2���q�0,gC?�4��`{� �=�n����Kd�?D�\Jn����E��_l�r��wSɚ�$�i��j�?�3�0'�E���֠�J.�2�����/�HW��l�b�9� 5���������J-K)V'�>.Gt۹�`?3�K~젢�y��9��Ŋ�O�/���OS�H�KYMZ�w�K�j�pE�CF�r�(���Ma�����^
�<����AB��T ��������$0�����/�"�}�5�)���K7ϋ�yE�£���{�[�0�e7��q?����`x������̦|��S�/��zLm7������fE:7H!�F��a����d�K�[���~P�2�V˶�CA��v%���Ii誛ϋ�$Ŗ�)	$��$B��娟��~��R�r��#�Er�ڧ/Q� ��G�hHo1����c^�0�+�APL�7BJS'G-oB�������T�j(�^L_�Ƭ�£�	Vs"}��˨,5~��<�%/%֡�48��h�A�"�a��.�+1����0�:F��L��Ud߫���װF瑰F���ɱ��l�3������oF��o�$6�s�p���CM�x��h��w�԰i�a�TQ��z�e_�L\�>m���	�gv�赏R�~|��GA���@��κ�)�y�?�6�6mߣq-�aS�U���>������"��_M�e�E=]]�şнU��,Ka0���	��!��n�S����#�p��	����_�HA�5jy�&�p,.�O�������mE���Iu:Ф��Ƥ�A�ȏ��:<Fd���0�@�����Q�;����^��tzB�+��q����S��?>U�j=�	]>������/S�`X���cx��?�1H5��ݡ��=��W\��ʨ���͕ޑi��0�l}aHkW\�p�3�k\[�_�^�j���IE��dQ�_�<N��x�"7GZ.¢(�2�!D
f�vB��=�!}pba���1����;�%��dd��C�i�4N���yT*y�k�I.d#X?�]R�Y=�����o� &�d<�OR9 g��F��}�Yx;��;Iv�,��X�~V�����L�ة_>- �����Ğ��y����ΐG�A?ƅ�f�E�������d
�_]���ba/x�D2T$B�~����H�%�w�ȧn���*y���z}��{�=�"�]�6���pnhZ�Hև��^�f�BpQh�K;�TB�Vx���:M����d���|�]|=�<6�l���ze���!���%'NKؚd�D<����;E��Av4���t�֖�0d����*�P�2����L�1���ڽ��M�a-�心�b�FC-v���~DJ��H�
�IQ�ܯ�W��F<����,��.	ڵ|�Q���Չ�W}C5�Y-_�������}���,�Il4?�^h�s�uڱQl�b�D�̔<�;=�.,Be�`�#�\ЉH&���p�6���7�)3T��믅���mc��F������p5j���i���z�)�!���{Q�G�6�K&� �� ^���jM����I�1�����'�7��G��\Z�l6��L��p0y��VXd��"����9����ɧK�ZB�S�eS���-�%�TlazG*�yJ�Z��Of���6j9BR�+��R����
 �|y��SP�.�ʝ�4-�O؜���V����{f�$���F�BixM�hi鸕a��B^����������g[9�1��d"��٬�&D�뮋���'\�w�b0�;�OӤ�,*�^���>��y}��;���kX��-kI��G�#oX�	E�����ߣ:!ْu[��'�|R�
}�g��#� %6¾!�>��M�_tC�h�ʦ���%/'��&�����l֥Is��D o_dO�`ģ)���o�Zh�IJ���������N��̹�GX�������j��@N�V��zB���Bo��CPn���Y��Ng�رM���~�׃�Ĉ�jS�[W oS#����%����ax����ڪ����a]��`_�C��YO(ӓ���\���ޑ0�����T�J?�6H���}]�v���|��o��W�����-��\E���ÿ�x�������G$�ɓ3���ނ��	�Z���"G]L����L^��/(�v������a�R��b��mC��U��H�!����H�!��*I��N�棷i8o��(l�PN�&f�[��_y`�v�8S��R��f��>���7]��G*K����(�h���h�׼Rͩ�J��E��v^��xJ }c�N���n�
^��J���ˏfIh?r�_��ј+:?GEݷMx���w}i)�{�9�o�d�ឞ�.���Y�\�|Ŵx��e]���\�ӯ�3+����er�ܣ�Tz�D�7�d۷�((n��ǣ�����?$��ć��N}�L�pt���_MGٛ����!��
�SDg#G�>��&��3���Hǟ�Lt�8/7H����A뛝��Qm�S������S,�-��������ߏuQ��؟�?���t�fS����"��΍��-b��7P�P��*e+��mBe�dq���`?�93m9įp�Xo�h�x��H�6f($~�ϋ�����?�:�t������t(x*M���+T�^�.�����7NK�L%����/\	ƨ(���xb����\�eu���7�����M�d*�.��I���+���?��I\5yT�]ǈ���;5�����~�����7n�p�"��c�a�+�V���ңr]U��U�1*7�4M�)��U�R���������N�����f�K�Wu��H����2�\T4ʍm�|�f�Q%��#w���x)!�h�+�
:2`U�Cc4�&��*:�i)%U"�'	:s]�t7\�q���ۭ���)JZN�c�ͥ�����'�<:�f�E�<�]���$���[�ʿ�d�3�]��Gߐ<�3��.�x�y��a��4�{��'Ȁ"b����\ߜ;�S�^Y^�r�d�=a�f`�L+o�-/Q�|sNϊ�ݝL kbH����MN�L�� <cϣ�.e_0�����;o��di4���>ږ�6�u_�|�ҍ&iα��*(Jv���t-��ӵ�Z��T�=c��"o��ݪ�8r5�?��sR-+>���ʯ�I���h��r�wS�]��+g{nܮ�=�h&tw(6��q�����̂�;�G�	�Z���;fK?�9.X���j��!
���jT=�Эb:)�);��o�O�u���M��X��� �3n�W��(W���֟�e���F�;=��Q=���8�{)��A�-�:��.��I����{��uO�	ޗ*y�)
yS�DbG�ݣ�8���V�/X��m�Y>"O��&��e�x�G�X�唯F%�)�^E�j�-:�<���� x�}����"�EZ[�R�
�kG&�$F��lze+��N�*���&�x����^?�� sq%q	<s.��M^G�)ɏk(�{��~�����HV�d�$�$���ݒ{��m�f\�^��#C�<<6�.������r>�2ZD�i�I�z3�����N!��3��m:BI7P�zL~\`ʄ�Q��?����E�����P�&���NY0�B�r���8U^ ��K%�Aq� �iW�Gx�ϯm$���d_ES��qd3�uKP?����I�6��SSӳ�)�Q�i4�.]�5y|�u���?���y3
kz�aK�^G���p�ϳ��PM& ����	P觓��Y|'�b8+t����7x �B�\���k��o�L�\q�r�ī��F0��=JW9p�l���`���f�ǵ���;H�q�}��e�a�x%G��Ej�y��cӁ��Ԟ�v�n�b���a�=�?�Ԣ%�2�?�90���~ ����	d���f�І��S��7���<�؏��{���i�A<g�*h÷<�dxT�>bYk�
��V�ƙ�\��,��\z�hq�GOk'�I�	�S��'߂�9۾09D�'��"�@iӟ���{h�<�_\l��@N��ѳH�㼿0".ۢ�y��Ά�N��^�^�|輰��3��'<_��j�V���K��[���q�O+�U"H�Ӹ���*y%�)���8��0vo3/[a9�#�̌��Y6���v1���y��N8i�K� �؀	��Q�t�1�iLR��pT��g�Xln�V�����Jt��L��K�������x6Wo �(Dx����V(N��X��	�s�Ajg$�к�E��# �Ìh磎��AH����u����/�RU�P��}�8)%�v�o��Us��@�(�Ơɽk���y�/�U�}��=��k�gm�J���NU4�\�\�y�}31%�j�
�}c� e5 $o}���O�S*���Nv�1��r��l���7b����+[U~� վ�-H ���Dw�̙�S��ř鷲4�����#w�l�����3Ѥ���q&��j5Y��2i�\��n��M�.�;L���Z��=#`�l#�e��z/�h�7HI���bh���y3��$�%ಓ癓KK���[y�6�Ӡ��g�6���
��-�ӈ�dq'eM.E#��֮��� �2RBKUk k������Tvn�o�8*`��z��~Y�ik���W�?z�)B)���㘡bW�mD�a�> ^���9e8嫶�l�<Y����{����hmLe�*�`'-#תĤ�o#�e���O/k��"%��W����\U݉ӈ�@J$��6
�s��G:xy=���PH�i���}/o�+^���v�u*���,Z�����}���kV��soU��^�̍_�[�i�#T����#�c���xr�c�s�|BV�r[|���$�P��/b�sv�`��PC����>/��u�����[D@�i��O̠^��$��~�T`�lR����)�t`Z_n�?�_%}S�m1��H|�|L��2+E��Qt\ɣd����%1-o^�Mde�����CK=b6C�����I�;o��2��{k(Z�1^z�|Wx��y�hGa�P�ʱ��*ye�WU���E�ä"J�r#(Y*Bz+��z���S��%��r��g�/L�:���GsU�m��ώ'=VIN{����݌p�v�$y�9�Ť��R�}��B��w<: ����E� ����k���7�-�U�����J
��x�o��@���*EԨu>�@�j!�+���c
�����|��q?B{�ہ1"�7a�/��)�>�Ni���X�~BLWOR�s!"���0໼�QRVN�u[F_���[�rƖ)ߜ��eI�k���X�Y�%������>�l�E�M����ݨϙ��%��Ր	�S5"|���f]j��-`L�?�����@J���:/���2�I��%��:�_��L@�������&�4�-?�����",&�����(���ĭ���\�H�V�<8��ݼs�ѧU��U����tXM:�HK�*D�i�wg=+s\$��ѵ��5�� n%�@Ի��z_w�z��\��)a��̜�mT�5��Q�}���y�G�TU�ĪLH?��!��CP� �R�(�ݼ �:�����+2;��f�50	����(=]���SV�CM�ǫ�ǂ}E*Г@3��k�d��0�y�d#��c�33�?��x<�����w��]�/4��(OA��ԋ������N�-=5���)U�J��yԕ��_�8���N��'���lY~�����zj�$05���l�˃�|�`����Ǔ�=���6�ܟM�`n0���bfAc�3I�!bXJo��jő70@	�譲�D7`
�<�i�ǹ�q���'���2����H,&��83���R�L`����l�na�/�(c����=��o�*�V�q�E�HoM�&CT�Y<"kt	�^.]�QZ�^�/[�t���.^�$�%4c+�SM����I��Ý�,�fx�'��{=ڑ����-��y�,g5�aQ��}�j:�h\��� �C�G��d��������N"���3eg������X#���9'fҼ�g^+�H�f	�շ�c��;������y/!�p(����L�b�"�EM�n�3�>Y2II@�D=t~x�$�t~uIG*�% ٤��%��m 91�4Ɓ�>h%UN����)��	��(*�w'��OmD�c++ϸ#e#�k}Ń W�|.	FR��I��9biS���f&?���P�㐅-�E|����PBv�^����M,��2�!^�a��&��#ٔ�Ԫ������[-�[��Bd�-��nb����L
�Z�c7,�36��M��3䔟�ڋ�=��\���6;=��]	x�Ғ��
ɕ`6UK�)�p.�N>}����7�}B���6��/i
� -��Ue�0�8�>�5��F*��G���ʗ�-�(�]6�G��?����:��y���~�����M�P]jbbM��ё"G2�ѯ��_�Z�9�F�h:��u�E��A��n�
�7g�g�[�s��x�y8y���ϟ��Sf�޶IY��v`R9��1>�z�/��K�Pէ�+v���yl��-�������V�j�;�6���:^�u-�[����Gd.�e����u�ҷ2��BܺxD��:�g��_<xN�V�z��P���}���f�r�*oDޑ#���7g������~9;�g�@ S�g�ܠ��C74�SN����Z���>g�����枿O~�� ����~�n�(6�,�O	�s�x�]����ԫf���R{};�*U���2']U��3�=D��q&��6qطv��ϖ^����A�q,�)�gA�q�q|&�����0���$K�Oywo�V7ŭS�r��Az���3������{�E�o�L���>�cd�����0��j��xj*�q��6����l�&��͹�Y�Xq��>���� c0�e7ke�^�kD]�X�Q�x���-��93�v�� �P9ߊ�z��\�n�{WrhK�LO�9�T�/�\���Z��%0��\�X&��C�h�'�j���w�oaT�^�ObZ�a�i�����;`K
T΄�o���y��0:�,��D��
��C5�,���@/%u���i��U��4����WK5�Y��oq�ܟ�?���;	!��%Xa��""��N�r&�1�x�}��R�ZE����N��4��ߕ�a����A������m�z�k���8]�ٻuMj��*����Ճ��+��}��+�s�޿�Eɯf��Ԝr��+����g~[������3���e�Y��v��������O��?�:�t�����ә(���V��_mBq���Gҝ"���~(��b����l��&�&d.��}L�V ���Pȟ��jq^��,Jhd��k�1��]�UV/2���L�?�\	'�����:.�pa'��Yi�t�@w���V��Ug�VOծ#�.��zHS���B{�vdb�#��U�E���7`е_��LR�TG`Q	�3���Im�+y����j��.��#G�y�ѣ����>�b��+��H��R<�Hx��㓫��G���q^���z"�]���k��7�9?�d~��f*+��}�^����\h��u8�rX�frJc�?J(���3q|��=3�58�e�n��i�ix�����;?N2�����	Q'������fMr	��Q'��aR����OC�m�6:)ޔ��{�]��Oy�u
X��w��pT\�K��ɽ������F����YLY�2�*ҟכ=������2+B�����t]�Ӟ(��G�M�n@ׄ?c0�p�0�������&�.�l]g$�cZd^��CvV���aKdTQ[�E��� O5X�&�ﱹ�k�$ܛ+)q���oz�b��E�������G��;g�O����c�z��hbȽqj�hL��_����\ݑ�&���$�lαW�N�jKuԐ_%?���痌�O�)�'����n��%���ȓW��`S/�B?iB�n.I�o��"S���MkQ�ي��؋jb �BVG�r��w�q����?��>�](\����$6�g+��� ���<���8/����[�s%ș�K�� ��yx�U�����a��֠�r��]�i+�?��ic�Ӕ鍦���@�a��=h�R�ɑl��-�����H �zi~ ��`=z��{dX�z��t��U�N�2���K��'w���M��?[��4�%!��v�c�Z5��mV��� |��V29(�k�� =-��pG�Т�l�-Y����F�m�{�D�Iv�$��O
���_���Yv��锨[���!�2!�d�2@����X>���	rx�o��5n��Z"Úz+�{~WGN��VK��:�~Wf؞m��#��>$��f��i>��_�O�G��N�Q;3���>��V�o�R�ޒC�qf�}�T�9�O���gl��C��Q�[44�$�����v�z��/� {���wc���3� ��cWx�p^��@X���Bv���z �e_�*����lp�U=":����傞$�|\T�F��i�^"��6`L�g��QQ�S,jdD�>����LFK���a�3 Z��^����DWްh��T��$2�t�(���ΕX�_%p4�����{�7aȚBq�S��L_�[@��{��� u�g.�s�k]J_�ۈR���ҍ�����&��ǋҵ78A8��m�oxH�Z��\�Mv�����&�V��x�$�ܶD�"���OBI��@�
�R���=:��9Q�{0��Iu�+Q�g�rw�[f6�櫊���L���[P:�5	���6��1������U�U^Ou���#��մ�`ٖ	�~�M���t�St�����~$��䝁AƊ�	1<Κz:	I�S&i�y���gu��t?pb�C�����Z�x�D +K��\����l ���mu-U�a6�hǵ8�Dm�%
W�� �'>�f��(�)e�d�C��Q��4LiD6���"�䭖eG��������س�{;�I>b��i���e��w	_O�0�8�ٵev�S��:�/ڶPP���r.��T�I�?X������޲�z{�������]��3���#.��l����3oE���k��s��ߑo�������\<�����~�z2���G�ɯ�P���e������I��hn�W< t�[m����j3�pX}�����_���ב�} ��b�m]*�a�������,g��@;����hn�ۚ��\>ƽ�*�PT��a�>,��<��.S�Pt�b%��y������L�'ku#�t�������h�Q�����'��f�����p.�����p�jji�l�-��댨E4�q��	�ۻ���u�c�}� &;�(�X́G���{ĺZ�m�����DTN,����O��9u�A����"A��غ��2�ӕa�{yp,}�q���*�$ցZ��&�;��W�\���VX���{w��q������e
�\��|<6������l�9*���k�:w����	��Zj
ZѐB��/L�^)p�"[��X�x)�jm=��U����T$�XyGy�nG�R�J\jq��ΰriO{���4�'��.�����W/.��h�N�*��Fni����O�t|	��g�.@"��o]V�F}KD�gP�;�Ų��b� 0ݪ�%�Dr�%l��y��[��D�M���2!/S#B���l�}NoLp��e��ih�h�Z�j&gdZ�x�[���:����^oF�uZTR+Q��Jz��k�FM��z" EH��hp"h���3ؕY���@��}��`2��E�8��~d��c��v�������&kf�����ŏo���-�]lx�	����x:Lqx��V��q�l�� �?5�m+p�S�@6P�l��{�%�\	�`���.���Q�p{�%���<X^$h}����O�R���1�䇾M=M��tkT	D�;��aśJ��q�Y�'� dB(��ˢ������G�IаH��
b�4�Ȳ�V-:�k<ًx�C0�`ِ��uf�*���P���d��m�z�z�(��A��˿���/%H�5E߽v������\�tY���-�-�D���'X�ͩ	�N�yW�����x���>���wQt�F��-���"�"��bTt�Jca�{q��Y�� ���� �v r�Ae�;^��E�+Ѩ7l�v�����g�2}����d�Ͷ�n�eG����e3���d2�)��fN��i�Gp.��p�be���NF��#�ڠ����uE��y`Ǻ��A���3���w�+���X���<\�qA{��Y�������#�"AhK���\������x�@��Z��7���u7YPw�D�D*�\��o�S����]wa�����g��lq;]܋�a�h�8f��������c�)H�2�>�?v8mjӯt����C�'�/�q��w��}"�|�]7g�¡����U:T�;z��>/X��V��^��[��a��BeT�7�D�((�,˚Բ4�ll��2~�t�S#(���41�4���<�住��E�U0�_���C�I����z8]�AuM�+P�*�a�q�ݮ�ʟ�v�l6��8�>��3bX轠��a!Y4E�@�L�NZ���5$�T3섿���"mG��x�j���H�?�/I�*�䎡󴲥���}鍙�.�m���Gȹ�u�\(2�?�� �*���$rN���lȯ�)~���/}�;��хĤ G�ʹ������b�0[��цB��+�2V��Zo���60m������(b��aH�l����Lȓ���)w����j�gu�X���:����C>���zH������	�G�?���|$�.ՠ�^~)���s��a���c����֥oi�ܓU�;�'DtP+���u:Y/n��gO~�����B�Q�)���oJ%)]�ҟ�_��XT]5<X(�bJ�PJ3�` �#-JH#) a �HwK� ]�Hˀ�t�tw�������>�Ȱ��w�{�{�sε���-$p�Þp�!#���Y��_Nze��*��&�^,�e�"��N?3i�ƈk�VP�����5��QRT�J�4����iv{݌1�Sc��x��g����B�-�I_���H��Ƚ�������q��!��$CdJoY�Y/�JR}�eK�;.s���2���0go��S���0>9i��j�3�ʨ���9i,�_o�")"�}f��z���_�3������$~<L 3'��4���5��� =��E�<�B8�һ���~;�͋��8�a��ࠅ��~�B�&�o6���4��L*x���'����(xr�O+��U�)c���ʝ7��)������|m>
�#ͨ�O^�cʃ���� 1���K˯��vđ��"��l��N1e�[*ߍ���Pc��YУ��HE#�VGX��R?k��]�2ht�A��C�I�j�ߢ>$��і���Fo�1���V�\��0b���C���0�-�.DA�0�'�Zf(�E'�Z)���2(�X�2�qZM|��7�4�*�8�c��0M5\�A��Y ���Q����|���p�Y۱(��>�&�ݟuA=��@���#`=�=y�\�#%H��Q)X{�0F��k��*���R0n�	�AZ� ��@Jx�K��,�� #F@.~Z� #�)=6�̬��6ݸ��,֯��?B�G ���E*�j���NL�ʚkn�<1�0V9�AЧ4T�^�.�|�/�L1�Nh;u�y��5�� �w�=54�;�8~��.<u��qz���&�`,�ں��m�i7e����	�{?9�m�(L�%Cz����a�$�H�����;��Ň.gjq�V&�����O7��$�/{�L))�~��<]�� L�9�7�I5;iskRt��*q�`�
���.}���M��H��T��-���߭!T�ä]���w����!a�w��i���;�FR�����63�݋�g���"�OIVt�<J��8�8w�?�'13�0��>n;2�;o8�"K�8L�.Y5]�B�^E��)�1ǝ8t�n�l��}�5�=M��,��qt��e�8�����Z��c�8j�0��'�Ÿ�3���_$��P���k��o�ᅷK�u�.^�m�������S�2�	#���"�q�ᑭR��X�tGQ��(兆i郙iC3cٙ�˖h�j�vK)}��"�gIf��V?,�@�������H_�����y�q-3y�&Ҍ��L*�����<r<��W��Z���=i���T#b��R�jZq�����&q��vO1z"�:���� Wf���j�ٔ#b�:\q ����"{�Ĥ�#BR'���Q��wE�&}�k��\��s�_���։��w�`Y6���B����<�xV�]m4��B�'5I�@�u��s� ��}��`4�#w]mR�f��2��X��qW��/7]���A�%8�F-���}r�� %�++�F�A�5�k $v�UŗĄ?x��y���2{ı>N)-K�		i}��i�9SO]���즪����	�x�����s�N�`e��|�B�e�̭7�����pj����1�߸��q�aT���Wh�Ž������.�hO<6���{ {����s�Q?%w�O1�]U,x��kN�M�^���-���F����O]_������Cws3c����͋��6�鲍Z����t,��O2z�qϙ����D�k�p�̯���.ת(��m�ՙ@o�̒P.�8׭�o�FJȌ����� � �{�#�&���m"�1sF^V�A<S��}{�w�������4n\�6b����L%N?�b ����*�f��NKj�홰EhdtJ�{&A�'�G�|���ݙ���������\��o�v؈����]%ZȦ�8��M�X��t���J���[�B#���j\�K��T�j��O#(ܭm����FmZ��w�XB��+,�]�HB�񭮐Ld�@��a�΁%�B�0�UJ�`R���"��_�[f�-Q��������#�}�qo��Y�F����q���3@'��^�v�a�#����R�tk�_)#��h�$�z�3�1_�����_ZPS�K�y/�����>�[��/n����C���� <�Z��[���j[��䩷:{Zl��%�.}w޲QpF�>.��S_�!��P�7 b�uF�D7TG�^�Hԯ�[4ng�	QH�.VץZ�Vׯ�T��<���~�d>l?/������͋o�wU\/��D�~���<{���Aj&2���Ԯ/q�Z�G�� ��Fu�yL˵Ms�/��D�)����7�3~�K��-o�.L�p%���P�h���n�����^X�^��ɚ�C%�0S�_D�)3�$�^=���ޖ�u�&�K������n�:l���h`��=>��t"g��p*�\� ٽ����.��l[G�2O5��ϥ\N�j%U�]B��ğ��w�JH�߱~�L܋�Q����onV��z[�$	��RR�q��!�2�A�\�s���M˵�N�ҖQ���9�=�W�JR>�\8|�_�[i� :�jlq�hs�
�>��6ݷ{�=��	�W�J�[Q�9uf:�w�w������r�m���r�Y5��� ����%hj_Ta�xM�\����@2�t�N�f)�9M��K%~r�?���l;�R7A�K�|��X ��L��7�%��������������~��t��D�HV�� �΂T��BW��-�;2�R2n��c�FB��G�f2�� }⮠���F�8#f�ǸmG��Z�[[������s{�e�3�]hE6/!�bI_4�xzo������.�Kw��L$%�#6|h9�r��{�뀣Sבj-Q��I�u����#d���]�vRvH���eQP�x&�rKb6~�W�A��ˍ��L�{T1��1E���1v�j~T��K�Jg낳��Q�$(�+��m�'C�(\�h�c����*u��5;����|��f�R�%\Jj�VE�w�%��/PfO ���∘��^)vH�`��0�t�E-P��Ia�ùZwZo�(1^;�h�Z���������ZM��B�zM�*5J���>|�j��{�ٷ.Lq i�K��8wب�oMKH�+�>�a����g��pfQߡ"�<��긃�����M-�پ��܎�
4�hO�d׌���VOƭO)C
Z����/�jP�:<,c��9��6T����Tz�ݶ b#֙+�5J����^�X�of�+�wI-d�`������%���f2�Z��)IW�&ŸS�~!<�>!y�as��?����~�r��
�f�`��9�3��*=�#���l�ӱn;����<�[�pnk$"�T��`Z�{=k����]VP��;��Q���#5�dޤ^!�#.9?}���$pȸ��/�be�HG'�,WW�t5�42�qGļ	U��ؓ� "¤�$�k��yB�������2�{֡;sϦP ��=?/��T�����%U���/��9#���qXFޅ2���-�^~����1g7���$���P\ʫ�R|���ϓs+�E�}�(�>�	~��fc�ש��r���_�0l:� 
M
�3w�kE��f��׸�[^��~����z�臭8b���[s���WukTġNH�e꛰)s,��>�����'%Zi_fl��ԥb)� ��R�y#(=�U��)i7�N���}vy�� ,�!� �f-5��zq���x˷�6wʭ�;K�A͠׎Pf���P3Q���_WI�D+>i�!��A	(�9U?�ڶc3K�c)�,�^q��3�)`��U�T�qӆ8�/�� K���K�ԍ9��|���7 �qw��j��Mm@̟HM��?����V�3����e#�����G���a�{(��� +B2�ɾHL��{�Ջ]!�@��*R��~���o�O
~��0dԯ��j*d�8Sx�����fӕ�Bۢ��2��$��|��B*�vͨ*�� ҉����@��kD���,BpՏAl �s�k����}ը�?|��*�MK��2�p��=�u��V��U�۾���؃�����U]OC��XJ��|7���S.��e��}������`�U�P�O���/������D#�x]Z������g���89����P˯������ H�B����Dd���i��h��T��GR]��)q��A������LE��tT��n�]cf�����9�b_z.( �!��^$V�]1������Սh�����Vǥ ��}g4�T�^J� ��s��s ��-"�3�$rZ}}������kZt'a2�KCD���Su�M����]O��"9�7P;=����gM<����H���>��7]1��e����%��3��L������[u���V'�l��[�łE�r�]�*߻�������Q��W-CR?�q��:� "�2G#��R�vk�;�'���Z5�ͺ�}�1?�n��If�����CX��w	��ޒe�3Q���	b�f��t'nZ�}.�B�WW�F�W@�kЭ�v�a���I�j5�Z5Z#�+:65�3u��l�&�!����p�^f&�@��G��\��d!�K����Ώ# �������Q�o���Zy��z��� �k�B�l�*���j�#Ul-l���PU�i}R��,��ѝ��<�7O�:��v_m[�V=T��36ì�A���?�#U� ��X�TG��>8mץ�4�B$�� ���e�o{��I���f��50���o�2�L����)E\Wbc�[Ƀ��R�gAP��쩵�0[���LLMT��.���q�Zٰ�ypt-�=n�E�M+���);�f<�����]&�۝AғUֵN~�g��sQD�.*H�o�$�^��-���{�սw��oJ�m=�:vk�h�ih��;���+_�
Y����+񿥰�n�ˋ��ȿA����m�nEHbpQ:w����XG^����^��X��&Y'�b��r�7B��c;�6¿�"L�G�g���5N��$�D��&|+i@���!��BJY�۷BM��?���e�^W��?쾛�:K��90��1���F�*D]��=X�88G� %�N��D��D��	٘��_m����2��@��?�\[�������,7�M��g��3�	L��T��+��ȁKQA���C`y�����s>���A�d'�7z`R��jF-���Iyx�(�j@\���A�GV0zftNÿ��]MJ�I�O�,�	�v=*�1��*?�*{�/�j�%-��z���2(��Ԝ_n�޾���^�d�]?�>+�~�l������d�8C�\�
�}��|��ons���υ�{W�d���t�7v(@�bc���=����,���	u�aS
��%�v@��h���x�(�B=M����}˙ܠ+ީ�=�u	Cè�4��7'�T��<Cdn���ݺ�*uS�]#o���DJ�4($�?	�}uBB$��eb���FH�����Fģ��?���:t'Lv
p�ӈ�V���������l�O�a�a��|v��eTȞp���a�!�S*���'m/A9E
�2��SqA���1�e���.��3��^�ٌ�����D��f}��t���7#��.�w��ˣ6]�� ��3<�+���������>��D��D�s��rץ��tnn�����;���}����z�+o�U�����/1��q�)A��Cϩ���S��㼑_�~>�=��2v�:9;M��?��iC�f߹
sD�5�Iz�ufz ��©��r�����uWfޮPQp�ҏKI�}�
6L,U+�G�"�;e���E�xg�n��<7~���/3���9R�j���V��RW[S�B��3�|��A��[뀠`EO�Ʌ�k����E�a/�ڞd{���9
�9�iw���
��������BB�^��=Γ�8��L^�mO&t�����i^�Xp;s�H�?c��[/C���̪_��c��RѳCo^�͑ q�4 %fS�/*C��hL1;u#�+��=�^��6x��������a����= �'�N@x	��؄@e6,�S�Ώ��̞M�πt8ᬹ�$���:���KZT�Ό�Ks%N	��D��A����se���&�UX��:�-.$O-y��0�UE�\���?��N*����#ذ���Y+��\ �"I9x�G��tr��=k�~=�;�'%�� W��/"��2p���n-4���N^�!��~������P�p��wN�=��o����0@�F2p��@5I�����d���L�S�^����{<�,II@�_xF�'̻2,cf�6���#)�4Bn����V�����;}�������������r���0��*��b�|�)���=>.h���tk�~Pdɬ�p굼�h��փ� ��F"���NA�_h�R�7aG��-yB/U7��W�i���|�'����O-�8JL���({HBg�n�]���kެ:�����rx�@NR.u�D5�{�;�8f�@f?�jvdϊ!!���ہ�MQ�x��宦kQ�{�K� �g���8��BϺ���F�Ύ&������:�ؗ�bu]�����UP&e��&�Nٸ��:��Ж������(ǎx� x��l�Aq�DL89����ǧ�,�֠�޷�A� ��`����<��D�ɕ6"�32����H)�J@=}�9K��-�ӗ���6x��-m�0T��9����>o�Ʉ����]f����fj���n}�����\+W���{S��tauV�B��T��ku�2�4`_+�y��.-�.��?�6����r�'MѼI�}�jgo�B�¼o9]�#�Bl��p�<��&����棐�~o�o@cI��?���w�jO�ݬ�t��i��w9���1�s,�)a�,厲Z�l�qs�9 v�[Zt�*wR��_�OmoO>���wÏkB��	򚆀��%U�m%"@#���Ƭ��]A��pP�fO��x���J�����>�cb��v{`g������L�-Q`k5(����T�R|+��C#·n[-,��//����:���8	c ��|so]偶w`Rb�7� ���ڎ��̩�c��1����k��wب���X�zcŗ#ʋwg�K*�����h@L�S��bp�S�� �B�~j��02���E�=�����X�6�JRw">���<���M���c�5��ߐ�����1��{P\ܚ9��:�T����������~��vZ�n�Ѡ�qK>�f��I�@$�K��q�z
45�����ٕ�W)�䥿Y��Մ������!��#홙� ��b���qՀ�O����@����q;�w��C��c]J��b�_�]?�ߓ�b{ �Sc���Y	��&�%��Nʘh� y��W�&j����{b��SL�K��I�o<��P�㤋}K�*��f��.�$��f����-�!��4Wć;}�pV��_���4���d"��w�;�<�0Һ�B��~��a{\Z������!E���A�����G�8d)�w�l���}b���M�p�6xT���Y�f�Lae_6��D\/p��ke�07}$�]�*�� %�rk���i�;�?0=- E�%޿����'h�>���,�#6��.��j/���L%� R�z�^���y+S$Xv03���oY�jέ�/*�焨w��.���#��� G��*����p@����C'}A}������j�h��4~?4�H�߭*��Uk�~,��\;�©~h�A(��O 2��46_��V�0���Kل�i��etG��.�`^����K7�=����_�ju%ǌڟ)^yEXe��s�`�G�Ǟtt�,�� |���)�:�6¯Xj����E��Bג�n���֚4_\@�!X�z �@р_g{��>�k�|�
A�s�E��a��C-|���PU;CC�y��J*e�A��e@���4�����"�` �ۀD-��4���~؄fP:��I��2
���>G�K4tfg�� ÷�u��8<P��{�t�:��wO�*Ao'2�1��5�1�f�/�t�I�{o}�lv�΀���q!H,��p�M�R�����`�8�-�K�
��������(�DF��f�^�&3��<1���J7J�f�������B�3�<0�7���j	&�
_	�N�;�	z	� �;�(Q�� �g������H��(0� tL��i��e����F��7Yٲذ���#�M���\yPU?��7��-i?�/�	���VEЎ_�纱\�
�;A���p�U��I�J����@�P
k�@~#τ�<��H�H'�R����/�!x#塺Ok�����ߝf4���UjmѠ. (�f8�j1�{�k�.+�v��Y����Z[R�r"D_��^O���5����L���A���!��ߝ�H;W T^*Zn��K�7S"/���aI�K�c��� T�qt��s�0�v  ��L�К&*Z��o�9AP.�'*EM�H-k��H�"���)屾�(� ��a�M*̛G�R�qK�����⅙phU�hSkW\Mɶ(T c����_�~;"A���� �b~|�Ms/Y�ͨ��	���b�}㻾�q��Z�m��
���5{��cx���_��L�;->%mn�)z�#�)��`�>�=9E���)��j����O��UZ0-����]����<Th,���U�B2!:{u�S@��|��#Brj���Z &25V��s��ى�ۯu�k�D�1�IIh���4�&��</TG�`X��Ч�QP�H�i� �0��C^����aJ��Z�ӗ��-���L�h�1���2ø`>v-���HMW��N���/���`� %I?QdЅl����3	Q;�F��}׳�E~�P e)Q�٧JD��1ڄ���&�&��W!EO�S���� v`M귐@� \\7{%��4c"m�6�U��t���U� M� 	���twt����c�yv�Z�x�dO?]�2J����Y<�H�y��:ʏ�Db�(m���?T��\ky��n}\����~�I*�z_ݚt��֏�]ݐC���������<�ռ��P+U�?�Z�	�����Q����>kޮU��:ӑl
�S���@�wI�⹘KXsK�xZ�>f�(��ӫ,�4����%��Lp����m�
 ��K�˴��9f�8����N�?Ha�Z���AIh�K���1�ʉG�03�:��R�xA�b�� �����Ɔo4��"g;+�z�r$���b���d�9��|)4�~��1�[�wkX
Dio����>NEq�j���m+~��p�S mfV����[��8s`��c�����<{��=��M�51Ѐ�&]���p�	�Pe]~#��NP���p:�?��#mقt~�����"6ʦ�^��\�a�����̑���7t�Cie���ø�g�}���d��}�kPն@!����c|E�	�[t���� ct}���qѠ;P����U�.$z�m�ݵ_�6�Z���`*@��s��3v�+N j�*�I�fa&��մ;�D&3���_�>�B29�?����`xW�����Q����31�J��H��,k�����1����v]�Biԉ��8�,���"=��{y���cv7t�P�V-�J��� w,C�Ԓן�Y`1Y�2�M�*������Tw��!}`Dn*��Ӌ��v+����P͏�0D��we���}g|��^C@��O^��5Z/{��Koڑ�4�=?�:�qƗ4�q;�pk�;L�1Wb�m�s�e�T���E�Z4(�	�:��&;$�yE�b�k�٥����1BΥ!-��Ѻ)�	pW��#P%�.0Θ���?{q�v˹�&�%��~���hu�D��wh��M��z�6��M/�;���vD�p)��X�=¶ZpFb�����������F2�`T�qy�2�%A'-��A��9��E9TX]��Krx{<j�B������s�ݙ{��A�2��m
���&�E����7��D���^� -X(�#�����u��r�j�G�����ONU�����2��L]�|�WI��-'J������v����9Rw7���>z ������!Y� uD�	���Ǫhhw�꧝=啐ɱNʆ���;f���=�X�2����Ќb�%n�z�җ���1�@�ye�Z������X7�ѿ*m�%_~̣�<@֡32��tkk��ru���~���@�p����z+��>{��>�i����$�P|�x8���P���\��Zr{M�i�[Ў�	�Խy�| O��q�s���T����|��U[Ec�y����If.�L�zr﬷��U���p魆^�t�jB-��nVY�T�_ĺQ�<�����|*�� �J�f۩Pau$�M���E}]�$��
Hu�!�#��ZE�&!�t�̰C�7�xc�&C����:���$$�W�^���C��	qF���q�"��nk���
;@�>k�/`o���֤�xA�a�;�d�lRK�k���q�=�>���]�J�j��$�#c����f����{r���)�&�1�ў����?�`_����(�}���|��|#�n�QN"���,+֭5�ܽ�;5�^ݍ"���(Y����Y�M�!sN;x���i�$3SA�d,J�c\��z�U+�ˍ���^�z�`��.g:�C%3�E��E�J|�H��v��!V�|��q~�m�4��(4`�W0X
°�=9��;P��M0�]�)qN��8W�uW<�Cn3c^�!�>~9L��#��iXV�]�J'����+ϓ
���.�CIi
���u���K�-A�k���.^sͭ���I�4b��$"���5��$4��d�T���`tj�m	�T�]�T��g��C��4����,����DӐZՊjF��!|	JY�h��6���앾�}�h]!E�A�V��Afu����;�`i�q=Ғ1�OZ�E�N*A�8GՔh2�L��[��hIRz�2ä���H��`W�&گ�{�3P+.� \#2�qXł>��� I����
D+�D�${��l��\�4�d�B���=�ҋ��;�����ټ9���:&6р0��#g_-DB�GO�G�3ȂQ�����u�R�y��T�B}p�Pu�����W��"�����6���)�ߔ�D6��NM����c革c&jJ�A,�� =�/o2�`�d�y�X������nИ$��y]�fR�t���R!���ϊ�N�E��_��F0Xt�]�"�+�a���K	��Z���r�ԃui
0�����sy;��/�Pv���z�+U9zz�E�y|W��V.�R1=*��z�&������C1է�9LW���r}K����������R�U����i�b��mUa��p�03��|w������xeMR݃X�g���"|���9Y�w�����-��'��ꀠ��^q���������P˚�Y�>.����
�S�*k-xw�x�N�-��@u;&d`�:��M�������t~.�{7���e�sͣ!N�?Tsv$�^�p��]�N��c���;��a����8VjpP�Ԕ��~O�z��P�����X�gU{��c%韊�$w�eS���H����Anq�LNP�l����
���B���aR�xb2w�,�tpL3G��N�N4]��?Z�
b �T3��y�Yhm}i2$έ�`���A���ƏX>	W��q��+|!$S7_A?�I�8|g�g�v\ ���2@߶��w��+���;��)��kh68mo����;�f�> �+� ��ȃ���#�m��b]ګ��mԩ�t��i甃4��9 ��o_����%��@���:��$,7�ߍ�Z�\�Oj��oW�;�{k&_Hr��G��v|� p�� ��iKgέ����R�D�_J?rOeL�R��z5�/Az�5��GJ��5	ST�A��cຎ�2=��RA�ُZ��Ha0ɇ0�����2�2Ĉfҭ�r�B���ݗ�E:�c�,X���ʍ�����S�]�qc�+`X����9����nYA̿���VtQ����;���ֶ-�_<���{�K��k�T����P�����.��-��Sz��[�1m�I\wvW�Gh�h䇱�u�k���]��l���ׄY������u_�_�0�-�}���]�c���U=��T0�Ԇ�W�	y�\]����E&�j�2�kԒ��&{��3��S�m����7��θ��Z��+�v��@sҶ'f和ҘG�;��:`�����mmK�h�A�
�W*vd"��,|���ë�C?��Zo!ϒ���\�˽l���O]��b�@�$y?:�Qs ���sKI��1��[]ך���MT����W�ʒ'�϶�bJ��U�~�$��(�aQb��Np:"�P2��X1y0O�3q�N6$�݋K:�P��UB���-��n-V��,URy�[m��8o䱕��w���<���`��K(ܧ}�$�yj(���]�j�[�\��h)ű+#���Y��>��s?��R)_@�6�tUf��P�N�ف̠�W[�`y���x�IXΑ&Z����E	��,�Ѧ�64��~��ddz��A�o�)=�5���.�;�D�,�"y�G���L��Bp�eӝ����sR���Z���eÒ��>�A���}���������8��X�6�muvߩve}�1�k�Y(D��ƛ�����8������\��^Bˌ�����S���"��t|}�ߖC�D�);L2�R���5m��<�r*�� ��yc��������|�|~�����@�9d��He�h�"+��`ׯAgu�PZʘ��J��o,*�]���l��!�I�H���zVd�����$?��E�Vg���G���1Z�K���.*�|N���U[JK,�E"���e���7��Uͬ����#����a��W��~71�eIM[z ��.(�Ŭ�=J���q i�s�Yu'�b��I�Y�������"��?�ΊŌb���`#���)�
E	40/ķ^��@�~�c��S��ʗ��Ii譛+)�[o�MJc�)��Q����I5�����{K>y��(�FZ4��"���VQ��z墵�Ij{䳡��F! ڋB����'B"��i5��QqCI$<��3t[]��(w)�|� 0��CW����n�ky��:��u=`�s��U�!�l'i�)]�f\�5O�S�GjO�6�����@�Ҁ�*Q�vb��x����1�j�����DNDk��&hAb�|��ݱ�qʢ��?�	�� �d~/^�>|D�(6t����i�|fã�+~�:	"r�7�,���ÔV�$h����/�.i�GWS^h�Y~�R��6[�/��P-2T��aXz�;�J)DҨ�cc8_`|�2(�^��N�{O�����ۉ$�]�ZQ���B�����F�ߤ���!r0����}�5�x\pҟ�2�ZĘѝ��Q����p�F	��#�ٿx�����Q�ߏ�������"T�I^�&0��@�;�/��>s'��\k�N����X�H�rA�eOQ�s���O�
�c/���؞��98�Ę{q�ڗ�TZ�|Ĥü���-����A5��;�	�n{��G���g>hm"��Ƞ���3y*�l�JrԲӷ����*ð1qɝX��s�̟�����hyR'i@5�����٤����;��E� Q�ɉ����~�
�G�LX������e�$�zz[;�@�-��冖��MW�c;�G�'��ʂ�� �!��ڐo�`8�����y��D_��S 2��.�L�-s%S/�ޭ]�D'��˗:�#;�gFM]������X,K��ή�0�x��'�[�=�q)1��q3��x&ĳ�؏��c�`��� -oF����
*�G�usjC�i����!ZYEy��A'����:zQ��bgG��!�9Lq��ԜE^��jc�ך��a��-�L��L��nY���e�� #P��?��}�z����I���Nɉ}��Mf2��{�,��+����Uo�p�����?���hAO+�G�e�39S�ª�]|9]��޲i2C-�&皛9ަ���D���f���w��K������T\O��z�wo2�$�=��1:��XM�|��Id�v/�� ��+E��ve�µ�E��dLjo�@���jw���� �b���4�ga��t���ڌ�����j�G��*=��2����纸�=%����$m)�<���8$%�a��,y��B�om-4��!@a��І�"X������c U����q-���,�jU�f�M���/�~n��+L{�"�3���%9�)�9�Dt���c�l���ff7EyA{&��Y|�sm���,k}ci����;3��{�k��s�a`F�ʾ���I6wyez͌3n�e�&\a�чpӟ��<�W|��z�sG]�ϡ�d]�'�"�p�>oNy�I+;i�v6f0�uiy����5zm	r�{�be�l{�qnӊ�[�	E�{����=�]�Q{|�BF�1N����;�<	~�Bumo%l?�(���7f.��RTw�fi�h�EL_nd3�o�t.�Sl2�7w_*�Ͱ\s1\&���<Xv�6������Q�k���H+c(tB�ہ��F���Y��k�;Άy9�6���6���A��pi]�,H �r���Af/��з?�Z{��#F����u�b�&a�Ś�ʓ49{w��D̊��$#��|�j�hU}$fݦ�x��{B�['NY���*|̈��6���RRĒ��'��kD�4������x�k���%4w����u�Y�5�o���	�w��
�� �Q$DI���$l��.VHe����#o�B7u�z��̂���K���VV��<���u�f��]�d�����D8/2��A��~V�M_���M��ܓ
��]�xQ6<X"l��L�v�ȣ����\��ga��\9�7x	�@������������K�n��c�����Mf��҇*-�zE5Yd m���ZMV�<�)��>l�4%�m�,I���jr�&�����+��/�GP�u��i�&(��<�g���1�q#�������UbP<��Z3$����bA+���v=o�
������k�+�)�;����
M\sL�����=��rM�Qx^{��&V�A�w�V�ɤ��`���,�2Q�ji��t�9�zJ��AЏ����W��e��mr'b��}���KlU�/���]�2�a �R���1F���,��=�҃h�qVg�Vf��:e<�h���l�DoӘ9v���ܐ$m�7�9FYS�^4�w�C.AL��>	��H�Kל��
��@��UXf��g��,��K+-� O0sE�u�a�t��Z�k!���xXCn����~�`!?:u���lr��E��хI�%��AC¯��'	u����b����^k
��y�4eh[��>�SkE��-xS!5�@���Ԝ���	6�5U�OZ]uk�V�G�Bcġ�@�/NQ�§k���%i/
��_�g�a���UT�	��YK��hi�����O�HfS
c���W�=��'��.�R���R��}n���#a�y�|��ߨ���C��[+?�<T2�Y���,����%q�G���OR�����26&�\�w�:�Sz���]�AzZ}!��M��>�]�1�!�7�L-%E�1�3#5���	g��Ԅ����
Ԥy�٫	����'%�d���+��@� �F�4���ɚ�ִ����iW@��� .��J3���Ƈ;e��❨��1�W	�ӧ�}3�j��6x�Q��� O ��"V��s��ur��D���g�1�	�����x׏���_������=����F��\��t"��@�8jx�zV�d�r*��5LfN%��<�`:-k%�u2R�ȳ�V<k�R�#�?�=�G���w��2�Y��ILU��l��b���a8`M�ffħ�V�!ge����.�|;ȩM�"��>)Q2a��n@�ꩇک���ox�F���Fʖk�P�`�3���-����6�>ؚ�r"�}�IF�"^�pY*���+p邤㦯
�#[D��_*�����ک����ҕ��GE7����s-��+�G�y��5��eTw��L��/�R)SE�JpR�F���y�3T9FI8�Ԛ���&��kS��J�_�yz�[�<�B=�V
�Rg� �}�
p�(�4H ���0�A�-�=����+&?���*^JG8�í����Ef��7�`}N�$p��#�m�Ʈ�P45�zi�3��������&���D�ݷ5'�X���Ҳ�g9Bjo���t�t�.J��Ed�H-ċ�8�S�o��饭e�ܜt$=<�̷	�n��� �W�]u��B�j��0�n�N�~0�D��Ɏ�
���E�m��0�K~N�-B�_��I.����C������؝�Kf��3�w��`1�R������X��'����w[�Jx�6�
_�%�nrB�u�]��U@	�5V�ٯ@�&p$#���^8)n��;1+�ft���%#�->h:��Pq�Ո���L���ys�G:yzh{}��~��/����[O�c5y�@ �Ἔ�mr���|��T�Q�%SǱ���J�&%�����
k�m�
��K����(�(����k"-�V����i,ջ�_raa#�zB��aW�m�e�vt�_4�c ����[�I�,j�m�Zr����*��,�LѰ�vX��"?�Di�����e������{4l�)+�b7�d����>�V��s֯e.�I
����R� �a+FA\�IT�0���Q����/�C.C2ĩ� ]h�m�դ�5�mP(�t9��*�D	���2IK��_SB/�����}TH��O�^^(��j�T��V�:����wxv$�jN��q���������aι�-�,���1-� ��R2�/ �� %�._x��9o`��o������������L0s���0*�u�TuF�ӝ�s�s+��^0���R���H���W|�B���)ߦ�����IPt�Y4Om�UC��2���#;�,�؄S���hY[S�]��n&�]�բ�s^#[�Dv�\��t愍�Ƭ������Ͳ�ٌ�P{�0����q�Ŋp������#^���~;���$*�8.Q�QsC暿�Qv�E��Fh��!-&�a��#BÐ�y��Da|�T9�.
n�'��;�M�!f��lRK�������+���V��D���C��d�blrz���&�}޹~Q�?��0���ىr�˽����LPM샪���E{��?�o����o-sel�m�}&5{�Br��v�n���ƟS	����@&AM��E����cs+���<��[(�����_Aϩ��r3�/���h�Mm{!�z��@���iF�!�&.X�=��{c�fA���P�ݼ|�r�
�)�?�����ڝ+"�g�[�T^��V^'H��`��3�X��8{��-���VT��Έi�Q�D���'��Y��;z��H��7���@U_F%�c3W��Hq�X�!�Q��J�%�z<�s��G���ȄI[ܝ��2���6
�=7]J|��sx�p���S�� ��m���u1=yeV\A=w(� �B��k��y1l4/�&�m3��WO�&�KMۄ#k���pR�Ʊ��q��@���:��sdSb�^Qr[�����FOs~�J�&����Iv���%�˩UB;%�d۾aE)y���V��9-Q!���A�]��Qugle�#��]�̪k��[�\I�.K�~h�E o0&u�lϳ@)�`�޺����`WS�����|GOc�s����%��<?�������gx��r7� *��+<P^��wL+eh�-���������WJ/[I_��c<H*s����{@�oG��$7�֏����q�A��:���H��̹)���W�C��2.���?>��O]�EPgv�M�=wǜ�<�j�<����A��
)��aaSr��SA��8s�� j�(���1^T��߬{u����EĖ�%�v1=�[I+)%�����ѿ3J]��k	��0̅���:�����V�%������?���_JV��4;`'_Ʒ�m!MF�(�o��T��d;��(6$8�u^kn�F�̅I�P�m��ı�S���t��RP)�co|��4�<M �0:�<�I���h�Ѡ_
�9w�!|��0/����Ʒ��"���ֲo���Hؑ�����������?��H(4�BBxdBiY�<�*��س�&ef��� {���M6���8�����=������u���k���}�[�,*{�Z�|~q�X��Y<F͔�ά(�w�#h�S:򝺹.��}�;eC��ÒD�S������3Uu�`,tϓ��*~Ak�)2�����<�,a���{� �]��Z�G��{	}����3�������=�m�;��_��n���ߦ����7�� �1vc�G%�6V<�y>��*�B�)f��щ�O�8o9��ľ1���ay� H��|‽�����^���	&�m,ˎ_J��?.}�����L�yWoɒ�n���0�!���e��xm��]�t�Qm�9�&_o��t��ɘWr3�7s ��KQ��?;�������?�wj;t��=�ۿߨ��&�C����P+��π����w����;)_6��>��QɌ�ز�͐-f4��}3���.b��r"2�3��i�;����)����^>����J�hY�����Wl�Ÿ���Y�Q�Q��vze��Z�4��\���鵾��t�WL�|x-���y��x�%+~�6^`��2������m��:ԘF��U3�a�S_c�)Y�8ҝ}���A?Sh�8�WĀ,����1`�;���x�#o�Ig���I��m����>�����VN����<���J2�xz����Է�+E
����ar��*����T+�x� ����ȶ��s�ک��/k��!m��4��1<�n�l�����gC; �̭DYN��������c^<�ΰ5�2>eت|�#�6ۊ�Mx�ݛ���5�;��{����#b��HNgN*��=�Nڒܵe7m)�mp��qU5{�
F!��(q
q뙧�%W��!���NR���2x����y��*��#���ø[u�zy�%n!��l�<�٥���甥��c��u#.�Ko����<w-k�p�*|/<�=�b���&��;#�1��R�ZVܑ}V���6PC�n5���Z�V���Fp}���1ލ���# \P��fUv�%�g��'~�	C�5�>��s�7�Qt��&�v�O�%���}�W,�I������}�0a�o�#�g[	��y�@�.{2��������+�Mg���6�z4�Nb�~����0>���Q�`�9v��f��[���%`��}��#�E�>���A���8S���,.`�R�){�ja�k~.U������e�: 60��7��,��­NgOj{5������o�zl��`�@��p���@ֺc��9��c�5�u�tz2�Ӱ���H�*�߱�|���T�kAl�QHn��if����Hp�<xΡ�����f!MZ��{XR�V?^p�717�T����gC��A�]�C�2f�/�)~77���ہOW]}���m�����"��_?yf	vݚ
(Cc�C5U��)��T���F���',.맊���}2)��~t�uQ4���2�x�[�����i�n5'��!R^]�6�D������i$@�@��W��G+	x����.e��q�"�c�b�Ys�jn5�5�g�}���~�^$B u���`q�
�����K�Z����Ǌ�`���Y�Eg���n{q�X���D��6�w��5@��;w�+·���^��9�41:�^�9�gϔ0�y�:���Děm�Wu���	��?���x}���X��y��3�d�a>�4�p�l\.̧��)P9��-�n�`�ڏ�@
��<BibB��T;��1~��#TP2G�+���A �A�~F��9G�j�h;~�竑?�\�q�:<���w/!�c�t�J����6�/����6�O�d�p�v�d>A`6��M�z�T�ʗ�HA�\T�7~���/�t��B���
s���H�,&�����c��` ���[iF",����j��|��3"R�.�ݫ�vU,�_��fu��l�z��������Ee��PBu�ۘn��2:�K��H��Q	ͯ����Z��}IP�;4	u��� ��`$o��,hsl�[,:m=��0���>����r�t�2ߐ�ӨT�����?)
���%؁0���"7I��)2(#��S#	����a�4��s��w �$����ǐ$�w@b�%�O�`w^��>���<H{	�%6MS�o���Lᑊ(��9~
����+	XU��n/ܵNg^i��M~z]#"��] Ĵ�������o��tQд�c�����K�ՆW:��x2�26Op�̗Y�{��ϫ�ٻJ�A\��(�'!d�5���<%3��k�L�b��k�aCS�.���s�W�ȼ[ �Lqu�n����rT^�/����Y�3tXZ]߼X��sH���5&�~7/u�g�*G=�'u��`yO��q.+~��ػ��n���@�P�痯����et�=^�.��l
���7��U��t-�@%���o|��ѹ   ����Nx0�M%.�9n�
���O�@�[�<��q\'�;R��].���{a��t �#��_[�������N�`��\���(���6��Zp���'Oe��S�m��s���I��BNo3 ta���*��ǥ�L�!w�|��ޟAԃ乮g�m��#��O�E����̀wN\gG..k���§s��E�!�6�U	�;�V죃�L-��]�x�Æ��S��]riR2F��K�+���7~�*ᯨ����<J�Z|�c���+m�v�E��µ�y��jB8���6�&�h%r�t�Q���XP�n9Β��q�C�m;��ih��&���#�~piz���Tn�K�+#S$Q(�����{,�|�����{ÿ7_��of���c�W1/W���u!�����˩���u��~�jk ��F彤��7/��vP�vm\�h�\}��gh5�3�)0" &&ֽ�����P4@`�����C��e����u_@�:t8D�)bN����q
��,�v����ԩ;o	T�
������� �v�r�}&���e��a� �N�i[��?�j=N>�Y3o�Y]=	�x����ZYW�"����F���f5`����9�2HiZMw�>��۩ofy�.'D�-��*s�*cJ�"!gC�l�9����6�`�s��x Y:Ww3̇��Y���C89�)iru�:7��s�-�;�#�l��r.X� Ƥ��v��w�ޤgg����[|�`ޭ�=.���O�keg/I�/��5�/����*6��He?g��~��E��(8�#��[츔9z<
�H:H=�h�	�Z��I%{]���}����e85=�|��������� �pA��\���ܧGxT��-���qJ�Bm�П���6b�m��� vq���	sʮ�0�*�GQ��0I깸�5��;����C�u����P�?�X�nn�����q
4��C ��̎v\"�=���zRz'Ϭ&��Rt���/zuH�ن8��'��q�1�ʬ�m;Y��^^m������&�XJ��~R���~+%��OV������2�̒�V�Y�VUޓ}C�^��k6�⺚�q�Ҫ�p`��Ew�κ��+�u�Wrp�)VZ�<}�7[��}ڟ�� ����J?�%�n2 w��0��
�lp�;{���uW��)��-��&���_��[���?z�P �vԨ,[�s�2^�Z)��ܛ��=�9������G��|�j���~����l�������'�_��Y�>��l�����5/=S�t��@PKi��lK��G-����Xg��^�JUE����D�� ɧ�wfp뮕J"�R?z�����S���c,�}�XN�8U����?��T�a������b��h�s��}&#/�x�`����͔om�7�	�V�O ���rd�K H��m�
�=y9k�uM6�B5߫T�&�c�Hҷ6���u�p�����$�n���� ��!S)bOb���.�C6�R#�����#e�?T.,V^���b�j�V��K���U��o'dC�ܢh�%u��̻�?���+4�˝	y=N�Oݰ��jn�C.�w�.g�*�Cm ���nF�L��5������]�ȶ��`t�������wд���| �̉@�N�ζ ��c0FQ���V��%�{HCN��"_�Ƨgi6bX���o��˗���.�W��Qs
���}\߳�hQ���y��2��;���P?r�G���kӁ� B��h	E3a�O��t��_��4�)��P�	h�lx�x�&�q-t"@��vהE*�9bO?̽�|9��i���n잍m�S����
OqC�=�]&k�7H]���3��,�3��6�����	!
�e�AYO��xei�-#7V���=���Ӱi���r-z/���8���C���t��5Kj5y��;	�2���N]O��M�|t�wL!�r	t��O;�n���(x���RqE��ʨ���Z���va�Z�>0	�8�g��ꦽ2cD_�t�f��qe3����<wv�v��2�g��U{&�aٟ#�I�#�5lj���z��g=$�O��w�������j�_7�6�E}O:6��4�����Wc�[v�]�s�nv�����NFMg��0�k�<�D^�h&i��ML������NC$�y�9ř��Oy�|d�3�2ڮ��:�K�7?Y �9lg��<xe��mS�*�����������;;�HGh'�]+�bE�G��Fθ����0��'j_�K����hՌ��L�Xn-�+L)>��*W��V, 3����a�y+e�{e,�ж�����,�G���|ꍜ,��v�1�л�U�q|B�'D��\����4,�"��\v�����HĮ���0���:��yp��bo	�q*'r�p�&��b�T�y�n��><e*]�g��?Ld�Y��.~�Ͱ>%&��7\L��a;rϋb-������������@m���A��#*@� �'\�F6w;��'^YU;�#EZ�_*u�\��5��m�Ƕ ���x"I���k��0�|��/.����("&�Gġ|Z��S�-�'���}^���г+S�+U�<@���lP�3O{v� �+�-A�"�Ń9XP��)��I�u�r��B�4P�n6�j-|��T���٬���F�s�����g+`���X�9w�kOhl/W��cUgps��V���'~�ޛ)W�4�\��\�v�T5�8]}/3�ɈK7_e��M�'�RJ(�\�Q��!��X1�9�(�������N�ʀza�����x$U�^��y��	_�<���́��)��f�s�Z?�F��j�{�58�z��:7��ٞ��@�Hw�}z���)��f��܆��d���n���MM���?cA��P�rj�g����N�_g㈶#v��6+)l)19�w��,zM\�^�0�:�+��	�Mr�|b����)�Q�CN���͉�r:	�>�& "�A��O;E�	$��_�)�+B���e�%�&�5��+Y�kn_����'�C���/BT�w�>��i[g�Y]e`���⢕0�*�v��z��[K�M󥇓;ۼl��O�\�y$#�������Ӫt��<!wd���cum�S"���[�J,����U�;����W�Hl���\I�;\^���kP���[����#��@5�<dL	��'{�J.A�ϐ��U��ި�G�ݺI�9cŧ���t���6和G������[�:O����p�sW��2�0�8����6���AQ�v�u���>����6���}v}��,�	��gj2���zlq^��:��yfM�#����Wm��ڑ���C�4�����Pg�����7�$����o'�`�k	�q6_Y��~�_C�����-K���)5r�0Q�n8�}�'�6����$�@O훆�?K?:���1s�ѐ�1���=8я#���n��_�d���럧�	���;��v·mڙǫ����@�5�%U%��t����焿%��&_6���0�k�>�͵����<m[��R�Q��ͪ�����]��\�B%�}�
����O�'�4�&���n��-��5�|i��p��rzK�:d
�	nƫW�d���[�PT�7_qL{��n��_��A`��[S��Y���)��)�����9����˩�1AUd����t�dj��,�r�����g��S��J�6�s�vb�|�R��r�j�\w����~�e�Cݫ���	��}�5ͷ����+#Y���n��0�W��O*ܩ�C�yQ���(��cG�]�}W_f�#����P�XLȺ	���hD-f�����M�5����v�4*�cQT0�W�l����_�u�����5+�������r�غ;���0�%�!+���v�����z��C��T�x5���L���2Pg*����3<'&���ٿ�X�TcZC������_��'��(�zO6�&��9%F=�jjM4T��	�Ƣ�g\g� �#5�O5-a�qF��ص1���u]Z=f}�Gyp�`g��.&�O�!{�˹�Un�p��5��`.U�g|r��i�xbL�r}�#�{�4ᜓo"![->�Z~5�'|�� �3{���p���'a�mA6�ٿ/��黊�!�o�#D8��
n��u�Y�b���>��7QܥK�H*+M=<L��	c�h���EB_9��R���N�c��E�|%{,�0��J����N�E�S�
�uf�� m��q��=�@�y|
2��2e�8�F��
�awV`�Sa�Q�`e����}�ѝn�|���`�-��W�;��%36^?��K7,���aL	.��=���P&5~�T���,���.��{#"��p�2OAO�
ޙ&�ւ�Ҩ��.'e��l�c�W[���kS���ңW,�_�9;xo��bt6���G�,�,�?6�ee\�>M.����U�te?��R(��h�Q�h8����I����"�6�*����
|��Nb{$�ճ���
�����7���JfW�E^U��/:��R۰u���wW����:���|��t��wu�%��JR6+�f��k�u�a��>����^#ٶ6g|�m�d�/������x�Ҙe��B�\�������Ұ�N�F�2��vڙ��Zn���_:/��}�T�n�F�;��O�ӊ�����ݳ��җ��o�rm��cvR!tk$��>nX9�Zn��V-z�y��~&O��l9Z���*���ٸ�6�4p�⼭�	���F������?��p�������D�����4/hUH�n��(6oP����0f���R-.���G��!�t��V���
F��-:����o���L&.\6������3Ig7��GS�f�K�4���Q��9+t��������r�,^�p?�X߻��J�iU7�ۇD��{jd��Q�"�,�$8��!�{ş?m;s���.��y��~g�Y\��c]�Q�S�|�y��7���}��\���An!��e����+�C�
y�q:փ_4�}��;Q�� ��l�>�S"4Pl��͓�e���A��j�*�wF��>3�_�wZ/ڂ�փ5Ҿ'(�,�ݏ%n��Z�Yg��ee�=���8G�7��$�����S֙�o\ ܀U_.�gA��#M�d:��_V���s�y|��u�8:����>�Y�_�
.��=�	Br#��xN�%B�H���5�f�"�,��-��̂l���Q�'�r���).�;<=��7/�^,�ώ6Z���>Cׂ�[^����b�	oA���b���1�M���+mA�sy��4��ь�FFI�>�rsI�|��*~u@�ꗙ��V8�ͦ��T�WPvUY*��{�-���53�����ָK��z�)~�|��U�4�Q��$2�%�ߴH׺d�m�~p�c}�]������5ka랡s����������ֽ�I��=&�Oբ�-jKW�m�<��>1�]�s�c�����b}���t���ѫp��˂�H�Jkd����f��jCm~b�!ٽ;{$�Fq���������i>_��v�\{���]��B�;���n {����kD��w�.(ԋ��Q-�_kЏ-ӱE#[?���1��e���v���cSdӵ��g�kfm��q&G��
���gtl�)fwQn��=��q֭ն����s`da�L�:�����"y�z���V%�϶M���3�s�M�.�>p��Q2��e/�ɭd���_U�k���R� ���d�0�Ddօ���x��O��*����c�����a0�P��=�U���.�a C7�[�7�O���`������1��LX�S�+Fn+�0��}*"ѣ�����zg��VU������Y��.����țk�T]��+}�9gB�}�:o@*�x�MOQyWq���N$e�	�&S�����^Ar��4%	f7=ۊ{	�g@D$nt��ϧ� ���$!!v��%�ٟa���j�g9�i�_����z��5�k��%^Ы-o"l��`BFf�ͩ��rq����ɯ�%�-�p.F�蠬ޕ���u�RG���C@�ݻ�q��G{!�,{-�����,]Ia�,ʘA�39c�ǘh��� ���4lt�dVڌ�k�ޙ �(S����"��R�.�[j�W���ẖ5��v�p��6����zr2�ټD$�Q�H�"��q��Lٟ���������z���E|���W���v�#����Y���u�G4[{7�=��u�����,�.���ܿ3�>�7.�-�q��jDˀ{;�lo?�=�?��t��	0��F)��=7��o�6�(;�w�cn�^���@V���f�+<�7�3ݞD��,J��+�6��wN�n0�	s9ݳ1d8�8��Cp�����@|%|����g1�ǌ�!4˭�pm�T{ǐO���8�jɹz���6w�,v@�pV��^B߳0��j[���� 	���bu��d�E��D�f��j�H#8�MK�d��<*fy�-���u��3�*��2���~=u�?ת��v�[�ݘ��X��8Y�cH,j�8Z�0x��$��I���֭\ �6�c�IuNR���B�w�O��7�J]=��P����l�/�ϐ����ߋcy�%?�#[�tH�e+��Ya�,�-Z�[����]`�f�ܯo����CF8�io�%	��G��Lp�}�c�]E��r��@J*�q{�����nho7ZG�����eQ]�RulIya��Mo��n�!�bN���1M�
��Y,-��k��w7,�;�X�B� ��^���=+f��IK��vC���/�O����r��С�>3�I����s���z�`�5z�5N7
�j��%�M��#��H�>�P����pvyړ�V��3T(.�� z���9��=?�,��'jգt ٴL'�	w=���+�.����ϭ��6<l��M�?���"l��5����8�'��ID;	�uj�[�T8}�(k��,�����`�a�̘H�LuX�H��gb��t'p��?r�]�4:��TF�A���)����*�y
Ȓ.���c<�ŵS��4��qPL87���T^�i�*�g����L��-z��W�0g�:&���QK��>�f������,�INg"��>�����-�w�lw�j���˼�m&j�����b�~hwh��A�����ئ�Y�qi�,�|�!� �4�X#��@"��E-w`��2`�e��d��pz�v�%p�mm��AY�m-�D��
S�?����e�E6�y*�w�m��}CD_�+*"����}�4�Ke�����0�s��DNS����~����k�k�Y�2g�9�#�~���+e 	hy�r��-p�;�J?$����L1�����=o��#|҃��J�<�`�����ݞ�b��S�D��?x�R�H]�ury	�7�q$+ nn��3mD�4��RCYq�"n�[��`��+�I��u�If��gB��z��t��y֩L�y;���}aI(]6 +[*�
��3����v�%����Ę4��M*�tn~s����g51�;C6;f���S~@s�Nw����Y�%&>���T�1 �T�6�wooFx��P���Iy�,�=��=ֻ��Y�*By�++�o�B��Tw6��Lf��-��h�N�U��Ƥ�-���(�}'#��
�.U�-G�k�� j��l�y�]>��t0��]�Jm�r��V��[���p{I�^�,�zo7d>y���ȭ���SB�+99((�v=��VL�~Y�e���?bк������6զ�׽�a��}9�פ��{�Kqv(���8a�ry�Y���&�-�!�BM�tXd�;�}�32��:��������
�dY\��J><�sb�����_a:{#SU}�2��B�Y@l�@��h*��#,�M�+Qӏ�A�����K�x�����V�BeRE�oc�q �*;�O:�e�&�����s�D(j���:�y&�K*�	�:�����"�j�� ���䑻_���[�8J����	�������o����M#C�!�?Y$�T�u?�2���4qO�9�[�E��yE����=LN��q�z��j��������5dxv�;�-�P��(��e���- Ɨ/D�9�-��
��p	�*����ȵ/w�T��F�';/�\�P��u��F�}�{{N����a��_�?q`�y�p�����.*�$�����V1�,�H��{Zm���Lϫb����?��]�K�L��$����8�����2T�����d�1H$�I��W�̈�؎��+�jDN|v1��Z���'Y�r�B����U�cu��tY����훁H� u8RV��mQ�c���\gvyvͶ$;�@��G�!snU�rb� ���ٹ;�A���#�T���Kuu�� ����d_��v���	3zN�hq���L)~�SP8��9M�8���D�\���UǶ�A(}��σ�z��-ͭƯs��KnJ�7�;N�M�)�����s��948 ���|�]Ei��a2#���F�P��� ���_�(���>M��D�!b,���~x������b�vl�ۧ5w�Z_8��^3/�7�H\Gwn���ji�Z^�!��Oш��p�Bx5�����Yp�_.e���+�Qm��^�Ύ��5r���%�x�dj��C�ô|��ژ��@�/�I���E'}];K\����� ����&x'L吊����q>�Ӕ�ꓥ}�������`���)�bƙ�o$|i5��Ԍw
8�'7�8ٷ���U��>'�q!��%/�	��¦�+��Ux,�@��@_[ט�{��&]�N�p���$<��,Yaz+<���l�ܠ��i���~��e�ĚF�m����R$ii(��+�[E��>��N���^w͸�s��M�|:�|������~Z����y��0c�#���V.�4d���d���<���$�@#O���l���/�lM��6���TY��O�������iǱ��=���1�F����������t�2�	�j`��Ѣ��Zv���՘���ɐ���wzM�F���˭Z?�?�[�r�:�08m�v�٥�7Z��ʘ�!\Ou���Wě1: ���1^5u]��N��Xf��M0O�>o�����l\^y#��jkԉ-���2�P��_��R�ZR٭���}��@���5�ܬj^r۝Y=>��[��K��"z���Zo��0B�^��O�%)*�x�wY�}���p�~�I�X
��g�u�D��ϟdm"N��8�������gGeG3�!�iy�Q���Z���\c����&� ���.�㧚����FB��Ӱ]�B��� �zAn�GĪ����z�#�h��!���qjXeQ�6g<��Am{�4���ݻ�&r�E�3���_�1S�Μ���<�+�5�Lj��|w!�\mf�JʥR��;�;'��R�Y�����+��0�)�{u�{A>*i	��g`+��/�^ώ8�S~>0r��j�_�K/x�Χ���qo�[�_�{�l����������N�i9��	)���0\(�<��q�/ɖ��-�
 *J0γ�aQm�W�!����8�;چm�����g#1~E#���� � ���^�4�FF�S�n�� ��d��D>R��ɻ���i��¤�I���M���� ����� �_�)2�`�|�_/��}�C�		�n$���^���'C�V�{�� �u���k�x��v��R���l��J����6:l�:��ek~#�Gr��ĸ3oY�c����%�-n\�eG����Պ>{�ޥ�x����0�q��W�p|���,S�n�.��ZsUd�p+��i�rε�]�yi�o�b���ɻ)��ڋ�Q"�V�|�E�v"�TB>	X�$�{�s3Zm��_͇��7�rGzd߸Nm�u���j�&�A��n�v�Ļ�IU�-Ў��x��8n�{V����/p���A&�3X����׹�7�nMW$��O�1@b5���v俬��Nϴ[�w�lbt	� ��UkA�Y$zl�*�Ru��nY�J�����}`���u��밠�JIٽ���Qwh@��%���d�]N���2�<Z��Vmo�{p���yx0ŧ`P숟'a���gZC�ș�1"y����{���'�q6���F��_�ArKoN����|�"�ϼ��F=T�;�������z+WsQ԰�AK�oY�5i��}�OE��5����'̱ŗs�����pL��O	'a��������SS(������Of�O'?�צ�@�@�ߪ���!Í\/�t&����%��������ǜ� ��N�מV��H�z�f֞�u��=�p=�	V�>+�⡒t��݋�ܠXH�4����7�C�+,��T���-<z�$��f ���}�FFY 5 wګ�T��}�s���WF�$�B��\�H�	1u�ęvԊJީ��*�U�4ɶϷ-D�C�*9�����H�)ۅŴ.juW��!�g���a��0�����X��ܼ4y�״���1D�P����r;�{���n��O<�㾫�� ��W�2{r�v�eO��ΎQO�n�T̝�����l�z4��D�STV'����Z��'�T��
�^�[��t��z�A�fE���C�0�T��Ԧ�����W$�{��b-�o��w~=��E-�Z}�	N��fXNn^`Q��m=�
`XI����܅c>Id��aO�b��j��˶�}�k6�����Es�}�Qܧ���ǫ2vp�g�SN9�c��J1kx�x�U+��%�w�������ڗa2�V#�H�}W�$���.��é�P���. d
����2Y�����냤Col}4c�2�ck�6���k5s�p(�7	`=q,�\W�����G<�����̂�Hk}��ʄW�\@�����T&��?���q!����]��iP�xe9Z�	���)n�+��=&r�V���a����?@5���'�(7�k���v�G�G�߻ތ�s�����yB8��Č�Rh`4CWX$����ٗ����#���~��o�>�)��M����3Ks�>S��ҁ��y`L�U��#�w&��#��/X��+٠
���G4d�+"P���q�cz��c�/��-�R��pu����1�f�ӈ��:KS�s���<G?)����"PP��W/�0=~�C��n��[z��M"ޔB�0�zc~Z����*�[��XT��o�"0L��>��ƀ��rZ;?_a[�h���F(xPo�ӽ{��(��~���\���͌��z�qz/�+�V�>��|�?Na�פ��5w����Y3�Ι��9I��l��c&������Q"��CP�|w{h*;�����]��Ƿ��f�Eˌ�ܶ��%��D"_I��l!�U=�8���e���`�U�t���`J���g��̀��T�0��#-=�=��NN�$���=z��都a)b�aw��$s�w /.���t�CՓfQm����G���	p����)B(Iu�+/�C��|��6���5�M޾�昃��P9L��'���5l�u�#T�˹^�����zZcզikt�^��~�^�.����_=_|Z�g&&q���5&}2=���5،y5���1��������[���ѱ����gOu|�=��$�3¼-X�3[�\���p%�8�z�q��.�,�b��q�\��	����@��'��������T񽭚9���Czt.-�}��J��$�=��nϺ�b���������((��d�Q����8��[f�BT^+r���9��WM��WN�s��j��<4D��>���M�Xm�%�!M���Z]x6}��q�|�3��]*YKN�����{�z%�{b�U�Ӡ����	]��t�R�ſ����^&5$�R�UH�S��y�h���bƝ����q��!#!��٢Bˆ$m3�jƞ�t`y�h����4R�Gq�(Z+������}4n���PL��^��-r�+�~��6m��a�9�,�拪����{b[*�[ː_Y��h��*����(U����+�zw�dCnu�y[Hb������@�|�6�Xϧ�G�T?|������zz���y�X��m�J`^���9_g�ڜ	w��zuS����V72����c@/5��L��U���PI���-�xj�3�L8�:��,��?:̛��;����%d��J���>�2�0�.*�b]�z���뙎���S�c�9�_�ց
6}W�;�0[UӶLb�WM���Qh�g��g�C0BƆ��C���85����!���]k��� ��e2��sA<�%Qw�\�.�7j�$���<8m�(��ٖL�6|0�jm�y��?\V�<�w�×A�^������m�����U���o��>�gQ5����_���c��C,}j8�~A8�*�����-9բMRj��	��Z'���(Qn·G$�m���>"��i���	���!�W��`}����T̯�are��_��ۦr����^���>�q:y8�-��_�,�@`s{m�k�xR�t�p��[y�ԋ`�*��\j����ݡ)�bL�2)�,��F-��`������#A6�m�S�S*@�)�%���bz�u��*؍�%G��;YLG涣���hK�����N�7�!�v?(���'�ߑ[%$�i���]w]�B�滽��n�JmS�=}~�Lc}m�2#� !8��*0�yF`x���Ƣ��h�O�o���H���#�y��\c������{�F�<���V�:���L� U��pr]�'!�P����1D�A�0��0ЦDt�)z�GB��V������==i�����6���vH�C#)]����ڋ�c��sC�EG���j��굑��T8e��%#������r�ވ2\ɡ$S}�\��e�0�(L"��	�Pel�m`w���Yҳ�w<ҫI�ț��ƹb=G���Y�����c������i�S���P�����lh�7�w.��wM�U�q|��*߈ʤ�9�1�t�N�MX��w�ޯ��f��XT�R�H�7�<m!)� aQ�/����|⨄���=��̐��x��e�/�%��[���Ǉ���t�H�}K�XL�^W;/{���op�N�\����M/�1�g�خ���u{o�3z�ѺD�)�yQ�C�}�z)�����$���g3ꤼ�4r�@r�V�Ma�W�'B9��@k���s�L���kHʥ��_P+MZC~^�b��rJ��`�vBJ�8BQ#��4��:�]OT���AW|s2=��vzw���Ƭ�Xi=����|w�����*l�8^���՝�@���/��V�Y����(��ӌOT�A����Jq[3�}���bf�F�K����M�Y�$��Z�s��R�hY�瀷[^��a؈Re;I��ō���%��r��V�ˇ`���٠Ā�R��za�u��)?�J{f�:O�mtJ��w�}B�;�9���1ڠ�R�;�B���2���+V}����C�4�FLr%Y�zi���{��da�b�q�%`r�
y�\=�Y]�'�Kű7F�^/�g�F���j�i�` =iN�ig�[u�;wz�7��M��Y�F��Q��{�/�q�Q�`�_! ��X���hc�X��n�+K"��Ď�i���|�W�(�hE�a�0嬇p����a
�`v��/��wR3t�O�>���"9����O�&��Z�F���`���X�x���� ]� �-��o'�a�lEª��.q�@A�#�v}?m�{T�U�.�{t��O��	�C�YU�@���{�X�͇aRR� x~�T"Fn���ޛG ֆJ��ۄ��2��8���t�$�:�����\R��*�)���o�&���d�1����=�_M���'��Q���8�+A+��l�~%F�y��-��ɇ���]�ӂa�N��h�J�|��]�oj4Wnؿ���k�3n�[I|;?�-K�R����l�@�I�5�N=c�'� H�	xu�?~_(��u�0�
�ZCH�!ږ�>��q0!�{R7/�a^_��e�Y���sO,S�,.��a$��|D�w�AB���IB(b�`�� ��/�.D��r��8�����Ywi�Ya�(!w�;a�$�sWҦ��\��2[�r^[�s�՜F�Ί����:��I�� Es%u�h�莳�'��=H���ڋ62_�i�^�Ƴ�۔�����+V5cy��]����e�}�S�&I��5s��Ǟnr����`��?i�b����)�����l��B���Ʌ��%�jS[{S�O�Hp����n��VI�'�s�q�y�'�q�����n��rI���C;��(-C�iGt������� ���
X�AM�ǜo���cݦ^s�m�"���=E�[F|
�`7?�c-vCk��m��ǯ�� �3T߳��L�_����s|+��o
u��
5��6 Ԏ��}'u$�X�6U$>�m�x��6��,vd�:R&?����MVr�ld2���ưR_s~���#P�ߺn"�|��d�*8=�<�| ��*yp����Õ�]�G�pA���Ci�M��O�i
��(4C�B�}��CPg}�O����a�f�i���z*���$wD ����%Z�u��`�iS�'*3�GreL�jmf?�<���05;�рo��(��O��|Ud+����c���<XC��]GG�RŴJ����� �:�vx ��1ކ
a�sBnye:���t����t��6u]����h ���䪷i�͇P�$BP���~�h��~�_22)�cі"�-���������gS_D��П=�����S�J�P������"��4��zM^$�Ì؀�	j'%�m�yL.��tP�Λ�&S��$T��Siܿ��F�)�hm�?���_	���кs�Q�2���j��.~(��'��]o�5z���D��]��.J�~h����
('�Iƣ���㞄���֘���^����n��7�c^z �B����q����%Ҙ�`��j��3�xr+��*�'W�Lh���P-6M��7�uߌMK��\��@��f8+e+�T;�'��# 3�V�
�����pp'�X���35�F����y�}<W	���v�MR;x��m:8���B��/�@Bf��g��7uYZj��� �@U��☘h;o��������B�J�c3��e����̑���֫��d�.v����
T�D����$��3��0O���D�8����WV���9|Uyg�P9�Uer���+!�"�!%�$%^'_�ؙ �|�PTI�?L����$IrF@���HD��2��%��dE�@��H��$�,�s2�����<���ݪ�ڲf��>}�/t�v��T��|�&��½?������WodZO8ۏ�w���|��q�X�s>4U�ھÈ�M�>�Y.3��E� �}�F�TO�ɯe��V���R�ݏn	�f|�a��n���篴B��]�\l_�Ѽ�x���c�e��
�U����%4ЎNjp5K�l��4ra�'Ӡ
U҄����Y�՟�����ɯ�W��RdTM�Y9۬Q�5�^�\��G�MjH��Q���ڟWP�����s"��q�U:��	��!.�ܲ�������L��妹��>�?e�$����a�9�$9�ۘ��>� 	�ӊ�ߌ
��ӧ��@�^�+���=����f�A��6-,�^�����E�9�Ė��'���NEؐߤ��p�S�s�_�JvZ�]ʦ�S�� �ս�_���VA�M9�� ��5�ΥH3�wS��H�>̖c���u��Tb��t�Ŵvs'>�/��drn�0@��F���� �1]�z-�Rv�		�<�|�E�P'�Y���N������q�VK���?� �@�=�6��b+H��9���g+0��Z�S�ߠ�Y���'#�~�����YXJP�]�5$�ZV�a��v'c�LEd�-����M���+P�6Q�P���jv���0��Γ9�6P7�߈�_y�G��6�}��+�tv$1f����#9�Iߍ��6p>r/=�]�9k�����\��� 1���'|��A���]�/��v�.�l��H�(��N>��s�5�_� ���O��l�+�<��V~�$�)8�qw/`����hSEs��7	\i�烥3��O��3�+�-mGD���i�R"%�⼳��h
��~��ZE����S�4�?9�Js��a��w�Z�zB(��9^:P��ݩ�l\�\5e�|�9>��0�op��<'�>�L�٨2���,|~ؿnw�'������t6C2=�����J�*�W�����z���K^�{K�ru_�xR:���/2�;Z %�w~!# (�LJץ:z]zF{�K�!�c�� g �{�\��E
��:)Zc;t`���<���ÿ��V�9ϳ��v��B�܌��W�l�p�jJ{✝M�e��Ю$�B�FƇ��F��K��0�'=_ԁ��O�� i�e������Ө�)������*�?iN]J/��2�B�G=���I��+�p���!s�_�M�ږ��}��)�S�
h��]���ݱ���"����0���;?N<9SZf�l`��%���\D��I���D��Aɥ	��,��^ݒ��%�L6��ծ����G(����tr�ט�iqG>��͚����a����SQ��K���fW����(�##����?�9`�F�"�Y[-�F�KZ�����s ��+��;(�k
+�K%)^�)ic���\<$�߽���5n|v���V(�K�@����:�&O�P��q�}���0��P���%s����������O:�i&���w�հR#�_u�]��7Y�黖��.?�{�'k���)���J�n�pq���`����E �����#��L���e�%Ʌ�[>��'��D��+�.^�����[I�0��"sP_��e���RZ n1�q"�]�w�o�/|�x{������&pU�:}D	Nwz����tKat �He`��1�n	��˰Պ��g_,F�NK��HA�x �Ć���q|���������?u�G�i�t29 ��&b@ӟ!D`_��+����~_�$e�����Y���{��m�\`/3.N~�*J��ߟ��d��:����9�d^���E@� �<V~Z�NM�Mx�P�F����_��<�����~�S��Mm�1M��*��S�x��^]�]j�s�(� ^ţk��^��-�?����ԣ���k��SE�2~4�B_�m(.�[�ܩF��FrF$-���/�J�G�Q�"�e���g&<'���&RJ۾I��]��*�(�Ӂ3�������l_։��V	m.��n'�y��#����M���{���6�~O�C�ꦌ"t7����y�~�}�}���ֳr���s����V*�Ñ�X��Vs�/l�WC����� �*���4���
�Lͪ��2_4��V�`y�
m�>�y��V�����S|���*���<�>G\IlK�,�MsO�b�6��Yr�A-ϵO߷�v���+]�)�E;�V�>�i4���������4W��o�BZ���}�����No�.�Ɛt�����^,���I3)]�N{[^�FJ�s�'�o[j�ɠ���H=�yΙ��:�tmQ���|�"r`7��s��:�%���g���5@a����[���j���7�O]�����;����.)�x�o�q7\(�4p��(c�R�D��]i��*�ʌ�J1Q,4�0��4+��w�}�dӿͥ�#����X�r{&S㳺����kiH<�I��������I��|E~�6��֝��`��ܕsq�C8�)\��'^��g�����nڡ�e�Y��fO|*��j�h�����A�$�{I�����2x�e�<e2xn��?��+��u�D��Yl�r�y��dԔ����z������̂�R=�Us�v
�䓩N��\��"[e�3���U�>U�_�o(h>��M��Ǿ�L~4�ϣ�v�EA�����˻�"�H�x���~�r�v�4�����r�q&�j�����9-��cbC�3���E����w���L�?����C�E��G��k��ף�~�W�a0_m�����Z/R�yg�{2�r<�Ϊ
�.l�;6'�R��Ouh!�6>���>ғV�rY_Ɵ,|�C�z�y��ot8�����U�9����[5�b�6�U�"C[�;X��r��_����U�dҫ�#u��S��+q���u�WQy��Gj~���)��1�����$-͎@s�e�KT��5�y��_[�]�;M��rg���^���	�
��xØ0�>�������пqs)�2���_y�b�_�+�X�ܴ7��U�s�$�?�0qk��W銮���Y:�r�h)/~�#o�;���<��h=a�����/��W�������dp�o'2<�a��;,���nu_[#XT�C��2zzf���L��⹤wڽD$�{'���!���X��Kӹ�ϳ�'r��::L���|amFֵZsJؽa�1�j�[�����g_����<q|�K{�TTاA:�leB���"<r��7`���+"��)�� ���O�ʕe>!����B�����ч#:�>[m}2G�q&�~O�-�O4Hf��S����_���� O�%��%�)����'���^c=dN���qn6�s.�$o�xjfQP�����'h���.~Z� �;����Ҕ�>�b��g¢C�v��ɘqZ,��f�B�]�����.�7�6�,�8М=Ɵ�t'�7G�vB���`7`{r����/Sτ�Tj|��"����u�Z�W��zpj��~�� n�hY)���A
���O86�J�ǕPyLa�x��`��?�@fw�]����d�Жc����������%#�+����W�ڢ�n�Ð�>���Ƶ0�ԝ^Ս���X���P���j�U�8]i�/��"�+MH8�4��KMݸG�����G�0�
鯓g��ܠ�g�!�w�/ڿ*U��/�v�Fv^xC�m�EZ����V[q8.Z��5�,�X,�s��_����f���"���΀��v��z:���D�ih���W�����#z��wQ>��<׸*9�݊F��nɅO��H8���d�;W����y�ONxs��r�������G���kwJ,����U�ΪY�
jT�!�
]�vZ���7/��u�yM� ��J���옺�ƁJǟEs��#�|�T:��3��S�s�Au������'\;<�a|����$!E��vl��t�w�Ls�F?Hw}.�E�3ް��8�|����?/�pdv��Or"�_%E�c o����(�����T^v�kY�U%Ӗc��x��-4D�ka��8+��I�W�.���a�k��%�Pr�5o~EmR|��^�522����4ϦT~Ou��x~uP��=dPHZ�����1k��3\�\��ׅH�G���|*���n1zW�+6�b*�˯U����(��!�x� tz�e{mu@0)��g@����}�n������ABu%C#0�N}������z�,�9�_�F�s�"����_&��?�M䈯.�=ffVg��/�3K��=�-�I|a]A-Fy}ΝM�v��t_u��E�'5f�|B��Ű��}�^��������!��au�{7<�����/���=�A4ސ� ���s���	[у"i���U��X�V!�fז�FyQJ�q���A�妶o�tAJ��.�b�;��MN"�EG��Fh�D�����Z[]��ԡ�����T�0M��+[�a[�����>9~��#��j �����]��Dp�o��?<���Կ��|�3��e�f?ܞ�ޕ��cAn�,;��r0�j�;�`]��~5.^�����\D�\ށ��)VE�H�Qp�rZ0��O�GTa��!��~��𧢮Q��zAZ$cӘ��HA^�YJ�Q��#��R�v��\�w��U�!5���7b��U�.*���Z�<�#�|,�X6Kǹ��J�%�vsR�:�V��`gCz��2�����^F}b3����HA)b'H���X]A���'���! �.Z���k�mИ�VIB�Q�A��v�̸�@_��9�1t�V�rV��8TLJ3���%�8<���w�MqNM齢�Lʊ�]�}NX~[�ʊ:���G������
2��Z�Ҷ��0^Aer�g���9�^$R��g!4K��Bza� ]�X��!9^�W���|�7�)O� �_(�~(6��.���r�����N�
t�X��G\�.�!Z@jj����~q��*�@kظ6sL7oj�,�C����F��GD��4d��*��xO�e�H�����9���Ֆ�g?�x��&U��/͢�-��.��3�qb��H
]5���=��q ���"��� ֵ���J�ԑ�����:�uB��{�m^��aĬ��pry�ɩ�ϭ|D2y1�߀�ʷ>��z�K�C�Z��!��g iq]�_!�IZc+�-֧�t��rӂv� ��4��i? ����дz��ݪ)9�XW�X�4Kݏ|�.L:��]m������	&�|��E�O�wY/׵��|:mb�"�|��9�|ע��DF�9���g~�Q6��߹�av�ET�Hs�sRy���/�,]r���X��F_kY���%B�2R7@T���:O�&�	>��x��6o~�:6 ����J_�9\5�/�����Z?��7�������'B��o�=y�1(~�+�+Q@�ꡩ�B^�%����r����Nu�T�\�VfJ��.�#��Vf�_Qx�E-�<�mˎe-ci�K�B,�egY}9lu�@��d>��lW�frV=�����)J�:��+��DJ�j�xXUGrF	��G6�@^�����qR<���T�#�<@��c�^{�G�k*�AV�-%#1^k���U[x��DI�SQ��G	Qn�\�~�ǂ�7c�Թ�mV��/�/�S�mO�S�O���'A�,�QĴV�oO�� i<�������{d�G�#%�eH_���h<����,F�MY��q�a�����GZ��YA}nB:"��2r4�?�yז9^X����p�
B��f��V�a���<6C-(^�i�0��>��mܭ�k����T��b�^9�]���i1��x�A��ϴguf	�����A����B���v$�{�9����3�Y���@�Vu���"����̜���%������1�����i� ���/���/�)�S���Ub�/BO�53�u�X	6ϾMK�+���r�I泋��dVg#��+*�]~˓���kL�h�[[��k�!��	_����I�� ,5H�C���'�Y���x�T; )+]�S}���e
�Cr?h�݌�p�������T�E[���W����� �2C��/9.�m��<'�/lH�k�P�c���ZX�O7Z���>\�-q�Z��Ч�j�c��_9�<�"ay.P��ysc�Xq:(�P]��W��d&������ i�n6 ��UA�H��4�*s�\Z���I�����W����V<ET̲rEI�0�T�욖�!�^P}�~����Q����諍D�D���|_�n^��f�@QQ�ޓ�}�uMs"9��|��Z�$k\�VX��o|0��>�x����ݧ�����C�#�vC�7�/�Q1�nw��z�P�};��P؞����pw*`ؐ"��ފ��ʛ_��MZ���& ���j\�e��Qw)"�c,,JC��3��!�A;]o�HU����i�|-���
B}S�"���Dq��C�J��C��u�ңUۼS~�����)��~��;i��R��i�x���������H�+ͭfK�w��w#�?�d�=�H�����7�����t�G����f=JG�R���Ƹ���}�8-��Ѯp À�b�� T�,Yݠ J	�����Ɋ2Xi��݃����ˋuw�H��1��a�:K��G{ES�{��Q��YF�֡L7y���&�d�S1��&r4�d%�
⤵�?��E���~vo�aM�ը[ z`���_@i����PR��В�y$�	0ʎ(z 6�A�䯣������Eh��Y��zޗ�*0y����p�����0�9m`��@0�?���Z&�!�T�W������*M��x�Y�P]�%?�n1nX�ʶn��#������J`�����Q�(���xJ��+���w���]�>��Ϯ�hf-(�����ڡj��M�/��h ���j��֧�?{��X�*����>X����2�{S:�UY���k\���`�@DO e^��czs[��l�YXw;Ϧ�+ܙY"����� L�щ������?܅G �@Y��q��BJ�E @��jv��q��${��>��M��g*\H`i���<`Ǭ�_����q�Y�~���I�8� 
-�ۃEo�z�u�����-��x
��r�J)���MJF��n;�w�~��7��O�Z���{���D6��s��� �k�hP��,/��y����j��Y��]�|Ȁ!*N� ��Ch��������nˀ���fc9V�4�K��L��ŬCD@��" ��yY�a�l��׵C��n��?�w=������t�D(%�e�ɔ�Y���9g��O�/����%�y���6?�S�`�a7^�+�f��G��9+\3U�2�䶕�a��$� ���0��9*���S�?|�=^��a���\/�q[�3�1{��ҋ��w7���X]}rv����]�MIRH�pq29:���B=n�{�J���} �*�r�����6h�������z�Υ���}c�YT`���YP���~�F�������M�B�v�Ole�J:u��M���'��������,��
]+j�H<������'y/�H+��M�t�'����`39 �c��	�ϒ^Dad�����;��c\q�Y�,����uj��z�)��)Ƌ�ߖ@7��;�bv��(�qg��T`�3a�jk?��Z�Z�so:��~�=�JU�s��}r�%�*Z�7iU����-�6 !����v��}pB��?� �z�j������kd��[��Ί�_�O��� 뱲���e��!;ǅ-���o�n�`�#�mG;]��lĸ˗���S�c�r�~�mGGD6���J��&���q�1����(�F9��mK^��$ +�>D Ex���!A�U�SWu��| ��)�����~�j�L�+�bL���4�S��_+���'J�G~Q������}�k��]�iֽvh���L�[� ���-� ��R޾��C,��5䬉�PE�����4�)J��{�q��J=�w C�b����Q�'��Hk0"�!�38�ޙ�;�o��>1�ġ��ò�������͙`����9�}zh�)֘�����ɕ�7AH� :�BX�6HNL@dD��_��m�P���Aa�WB(%���$�U�)pO}���^٩��h��a��c$�)���Ê�<cu�J Mj��6��=�Y^{���Kx8������L��WW2~����+^fW42m{���)�
��!){3ꮰ���"��'�[�o���=����HAXmE���f�J����W*����T��9WP��O�$�fA�d�����o=�d�5���fѼ�v�e����|���G�;+�r�.gj�b�7��Z��;�5]�b�'Y�DQS����4+��Eu�"B{����D�!���Ԥ���3�1k�CTIF~E�o.>�JFgpҲ�DQ�(��Ȧ��qa�1�J��%�'�~�X� Qv�J1֞���c�����X�&U�Q-�C3����Bxo+�2���mx���z;��"~� %��.>3.��,�R��o��mo�2_s�)�Q����*}���3�ps?Z�K8���jH�-ֲ�k�[��_[k��7x�����I�ń���O3�I��]5Q[��Σ1�ŀ��ή�`Y�ϐ���4`�Dj�h'���̾�=Yf�(EKMm��;�  �E�W������?L{��X崄�Y�.X�B���l����X�w�_�;��A�W}�vNZ�b���!��~�9�d3��9���u�����E"���?7O�(�]��%�+�/��pc��~�&�m����UK�*"��C���eR�OnIܾ���>CG�B#�
����E�������,6��g`�	A$>�]o�*>��O�'�:à1���z��������#x�w���R3��X�Cf�
�;=R��:�,��vc�������t wl�RP��it���2��4�<a$񐆥��&�Q�.��^�8?��?�r��qp�����d�+/Z�(��J��8�*��P�k=
	� �.��_���F��~��_�Gr
�͌f`qҝm��N$a�k�Q�@6%����s�d/��R�ܙ�*��0'�cm��!-/S����%��~��:ؗ�bzSK�tk#!�K(�Tm�t�xgs9��n���u����eÓc\��A�l���̛#{?���G�t���O��F����a S ]�������8�%d�xl��K<hn�}��{4��e�R�����Ch�����X@��,P��4��?������'�rT��v2��� z������r$_�����Tz�q�s� ���]�O<�&�"3�Q��c~� �t������7}�y�P>Lf����F��h$L�	�����SQ�{�0t�,pI�ϯ���܆�rt�k@� p�mH��8����q�|��@�Xy�jw�zO��檶HZ�Gt靶X���S}b�[�q�ւ��}G��g�$��u:�%��8;��q���V�N!���|�|6F�D��x��t
����I	7�w|��^B�|����k��8����_;<�<싟�2�8B��	*Ϟ]X�%h���9�8y߉�j5S5��U�>�4]���ɸ��X�⿘P�v��g��	;��>|u���H�cd7�庡g2w6� ���#����d�4��M2Y��އvv��P�?�s`䣱�9PO4r�]h�x�)M~yy�45I�ݢ<��ؕV�L1�H��tz��4b1�V�Q�d�Y7��gG�U�-���lf��7�^7G3�c _r�`�o0���@Y���3;U�uC9m��]Ɋ:iB�������P�
3�c�c����#=qR�; )�d:� �x�R||_�������Z#$�&��n_����Z^.���W�K�OH�@���uw��@�)6ٜ�I%Z��.�h���7��]�K�ŤG(�.������2Oz���e�.|]�HF> �	�/�1"��b���T�8(4��DW�{��Ԃ+��ĂQ*Q�.�R�18�P F͡96EY�Qd���)�F�+ͬ����Ǆ6Zr��CabS#�IPu�l�-4$B�L��qt=�ncRr���	q�Y  x���?�
���C�����ۙ��&tڽ�#/`��z��_-���19ux�>"��/*����r�]�H�
�bR���VYbh���l�Ȼ�HNn��Y
�w�2sz�p����
�m�rk+7��f��s�r��خ�SǜL��2�c����Ρ�w.:D��Ϣ��{Q'�_k
�G��#���v�O�nSJ>�`��CN)�"J�!�����P�i�OK0R�M�J �M ���5e��;����o~X����Ǆ<����ҿde�s�QO�n��У^�y�ש8k�U>�8#`��$��*v����ȇ�DNH�
R��9QJ�%�t	~Upk��{o�@�C� )/�	�d��ydZv� X^ۖW>�x�D���Z#fE��� �@�9A�ڛapW(7�!ќ�S��g��eG��j�{�
e��GL��v�$��S�!����Ղ�?�g�#U��sy�Fs�S�W�㖢��%#*_V�ү�A �c�ذ;]}�!�y&���Q �t�u'���կ{he�;��L|��B|�v������4�W���P�������ԏ.���ĺϝ5$$]6�l���,Z&��%���H�4�\��sT�y�D~l�i��Z�����1>��G�#�.ꥤ���L�jav���������~E��c*k�?���=�%z;3�PX��y�H촣�"<HzMV���z���\�Ò�/�lS8PJ� �t�t�7��ꎕ���3�C
��"(�g�.° ρ�r���&:�I[�t�����U��)"����UY�Kb�MSxOx�����X�{4�g@.艛�_�`��z<d�f�?f���6�}a�J�9"g4������$�k�́�ꪊK�t��,�`�B��!`�.��������mE���$R���O{ j�q��[�	�B�£�!�]U;�	�!�?�I��8�����b��|��(�[ŉ��[���n�w4��������wM%�{�W8��-��CJ�cV�7T��\�e���X���i�QEz�`��?$>���? ��C?0�䧊�7�1��֭�遷=��J�1�)��]���Xv����տ���H��p����w0>�À��= *]԰��,�(��p���4]��@�K�������!W2[�b�0A�O^��߆�>����Ÿ*�%,��q#��VgU�ȻE���c $���;CU�I�����ߗԡ2��3A�R�����,��n��}֩B�zL=���R,�~�@.8�_�on���˹�)������6$u�~"�Kj����зU�l��������:#��b���W�
��\��TI�X��e�kI.ɯ�����Id��?F2ɀw�ؘ{����0�se=}S2¹��]�,�n�����h- �Q��|F������U=�_T44)�����6j��%z�8��/b��rm�)ޱy!�����K���0
8~v��
��J`�l�gf2��f�F�#H�Ph��oKV76�jZ%#1O�ഉ���7��Uᗚ�T�eP#�JUdx�V��AS�#�VaVU��F�!���G���k ��'߸�h B<|�O��w3��4y��.��N�T��I�J���G9|��Q]���З�{�L���u���8��?��=�\�O^�!�(��s���ƯV��"�.�K��x�W�&8��`臑�3���<%,�������@O�^-B�*��[�=l�\ؓ�fRV2�/�k��k���S!q&�fM�-�}Ӻʯ6'�]os����8��[���n)�'�a?�$Q(�|MZM�H�+�2�Z�6h�nI��q��,%�$�7r �N�� -@"�"h������8,�
3�!�e�E�Y�����L1ˎ�6�I��a	C�/�sV'A�}ٱ0�O0�گ�{����~��b��G�"oi�lEf�H��
+��~W����N�f.P%��T�o�b��L��F�I�vv�o�!5�Hc�IԚI�Bd]:_�I�W��A]FQR40�F���|�HH5��o���꒍
��`~�U�5j�}64Jp������k3��6R��������L�� %v^wj���������{�m���)���Ε`��xƀ�8y�C=jb�
K�\�V%�<�)V��5����@ۇ�0�=|�m�����ܞ?��!p�&�D��<��N�,N!d����X}��k4��;n�O�.&|9�SM4�L��%�"%j9�t��T��Le����7d�����9/>#�*j7H�y����w���߁/���>�W�8���L�d��4�~[�h`B��S��M�.�9o^�;���)�3����f�̞.e�(��7��#�j�2�onT�Δ[�w�b��)��?4�*zz=��M:�1V���
�u��i$U�?���o�%�/�;n� ���Z�⭎<7��;����p㥿5!�G�&X&��vl��E�$
֋d�*��%��bY��H xs#������>�g���s־.�%z$���-h����c��/��E5PW��_y��x��5�?�g,��Żt����;/���?hR���c��	_��������-~F@����k��Ա��*\K��|D��" b3i�`r����:oZ�t��񕴽��BHV�o��i����C/'�_�ypo��������T ��m[.�܄sZ��
��G�`;����$;W�'�WP�����7�2���.h25`��H.T!���M�~��3ɢ�N�o����0m�5�'@�+E�Zj̹�m�������L��π��:���Ύ\λ��������/)4
�ce5ͬ�|P�^��:ar���ys�:�HџZ�� c��f>�w���,��T^�u�z窩W���*"$$�B����E+4�^��.L-p�nE@�����>�e0u��� �1��~���(���ul?y�깻+ώvS�>m �C�<c�����kZ�$������o�y�B����U���|�m����������>|�u&�9l��M��G�eL(BP�u�3Q,Dޓ�z�ji3Z�����R�]3��A��w��Z�	�_`e# j;eû��*�S��c�w<�Qݗ�S�6�6FW%�V�����/؞"�rd���I�,���mR��;ԯ�O����[�
__�8�x�'���b��f���0m��@���`���`�ܔ��.��5�7�XoPN��/�h���L���bm�JI��5�ݐ�̬Pl�|Xn�O�.�]������:+>��+o���u'���v��!���
�a�@Nn\�%2",+��1��1?��^ B��ia�q�P�J���)O(�T���!6��׍�F��e����&�>�Bӿ<� �-�ug��ē��M!	�!N�β�'o���$��k��'M�0�U?%�J�J�&�
�Z�!N{^�HY
��V���m^�Mu����l�%�w��gw��T�oߎ7ɯ.�Ф�h�5��G�)�òxVoDɌ�u�h'Q�����
�+wc��h�(	y��Aw�7uΧ4���6����hH�o��j11�$
���Y��8���g�Pp�o|C/-9@���DI�u����B����]kH�I+��#����KX��E��Y����B���
�z]��J��ao6<�Va�c=�h�rZ��m]��]�M�hj��Lh��n�D���!#S�Z��Ϲ����=B��%��-�{�
�'_	���T�qfR�}35x)�f�ڭՕz�#6��~���#Be�k�ބ>/_�[ �iM"�A����S�)���AG�6�~�a�"�HO���� �Ge��E����V���Ti�2�:�04e|C|����Z	�0�E^M���&�6�E�&!z9QĔ��,�/qrY�?|]U�0B�;�4٘���C.��b���&�`�$����]ʍ?��i��Js��&-yP����(}�I�y��m�e��6�6�|U�4��CITْ�S `���8�r���9X�~�5�P;���l��RK�����Z�T�O�j����M��,�;S�"{7��g��5�ߌ�8J��T��4.hÖ�s��*�K��m�����._"E�Q�PK��O/��9�(K-?�s��S�w2 d,}rVgWd�0z�7 �O�ɐ�,_��"�e�Z�:7� i����e���� �QS� !��@��h-27>/9i�]/�He�|�aZ�� g��@7M��O�k|�����;7���ٛ����y]��{�yP�H���.k\����@Aw�U�?r�|/q*?ߞ�KD ���n۔���\�kb��"k����Ս�w*�}��~1�f�����a��4ٹ��f҇���m�ײ�o*;�4��������*LF�I�h�Y��Tc���*��$�d��M�#8?��+��W�H�K���� O�6�p��{��<��0��*^n��#�����#m�m]�d�ְ��_��|�1g8r�����y_E���.i���~R�$�./\}{E��R�Q��ԙe��ߧX\�S��Җ�
U�ݖ�PQɏ�j��l�i�L�x��Z?�Ç��s�}�~�5�O��Ώu�ߝ�"�kɎ=���;����O�c�'�<��g;W�'�I'r�)`��P��b(#MȂs��[k���{L�۪��{��X�9�uba%��^���!��7D��(��ȥ �b����M���+M�Vm���G阆�]�y��Y�6�����< ��O��*��R�Oћ����l���Z��Q�șE��W7�{�s�i�?g�a�cD�y����cYH�Tn8@�����O8�L���i5[<�5��Ic�/�33.G4�7(_%E��^ dgP��Zx^�s#Я(5��^��ԦQ6�Ж��� ��سۺ67N!C�����<�z��W���t-Oy��.P8�>�������TC���KGg�������j3 ������F.���\�L�'�*W&��F����Z)�.�aiCO-.�[=��a�'w�I�7�hW�(��ض~#�8:��yAc1�a�֞�@ɟ���>}�FLAV�u�܅7	�nP ������/����"Z�ߵD��?��Hg8��y*i:棺d�^!\LzYQ��Ko��p�!�ՠb�%�B���-z�typ{�Z#�u��-;�i�\��H
a7|���� "��!k�؞����Bcɲ/SV>��0�y�n�Kpgif���?c~Bћ;9�9�1wL�Z��-�vT��z�����=Y"?��`}����sӱ��ؒ�k�'�nV=`����=�=Q؝v��I<���u�����K��vlOtr17���逎4���0�u=��=><f��"��Vn��|��(�a���f�i!r;"���s�ƺy��� �͝����u�����v��?��v�8N ��V�v$����?6C�����r���a�aY��r����q���z3�W��r8/-���<'�h���/]�ߐ`���_$m�T�)?T�T{O��-�ft�~L��S�gͷ��c�����0�]���,���d�K�I0y��`0G����X�\��Eu��΅��ݒ��U�
���ߘ�F��Te�a��V�`Ma���s쫘�	���Oa�����7��[���� �o�/z�}�
�����Ȇg)��4�m�i�'�~�_د�㣔�1��A����;7��������?����]<��S���BҘ�y�»w�>/�9)��޷Zfb~l�H��TO���E�E<�'��6��Z�	<�@�nq�On�t����fUMq�7�7{���V���V1�c�C'%��3�σ�#Sָ�C� ����i��i�����ȋ-�WVW:�Ꞑg�C�O6+/v��p[�f!�,�G���d�0t�,˦�D��U���M�n�i�ֆd�v�Vc���k��l���$�b*�W����+ۦ1^no6��O�l�-���c�M���5��xX�Lc/��O6M�f���{�W�Q��r�xu����!u��O~?���'��;U��n�b?Aq����)rm�%g��f��D��P�T�]n|����]����C����,55�[��wM%����k؊ku�7���C���:����z��K@�B:�w��N"e�b'Lܷ2�z����p�J��j%{?�� �n��x#K��������5�m|��̥�0WD鼧q�g��(�;>���=V��)J0ve8^Y����[�?�˒k�Ur!�O^w���w��8z��G��l��'���蒹�'Q
�j�V$���������Q�0X�~ܤ��<�;::�A�5����������� ���6~���v��X���]rW����g�܀�m�s�x��!gn�i������1]t,[op;�T�^Ψ|:���#��@?�w��-��jhi��5�C�x��;�i2/��i�������V+�Zz��M���evuqC��#F=� 2�*�ha��]�����t��[ ��c���[���w_hL���L����pG����%�p�д�:h�w��ۺ�(�-)�̪n���0�^�F��/ox�d�U�}n��`gf�hSx,�,�����޻~�2f߰%�cR�/�����P�Pܘ�:3nE��e�� k9��i4�͏z�P���#�봩��-�o.�c{�M� ,�ѹ,c�~Ǵ���2���gC����"�����Z�oG۱W~ú��y � G�fQ�JO���wbN>?�J��2��ֽS$M� t���Sv��:�rΙ��|��a�)4�2aPƛ�:*c ��uwl�@�C��Z��50�z��i8��"��9	:\�:�L\$���w!����꟧���[ G?�����Ŷ��f}������'�y��Y��� }qҽ	�����k��>јM.h?��}t�G@˃,���"	����P;�9�>E�U��Q��J��k[���*J�R7�����.++,��8h��_[��b��r5OAG�`�=�̾q��ԛ�p��xzoaw��ο����i����� ��_�����;��>4ү'�p��Ϸ����]6�VTk|�����[Lg�W��Ph�W�cЍo�$|�Pŋ�7\��Xw�pA�t� �+�p��?�v����A���W�A2���nn�iw��+ ��H�����M�'>n�l�1н��9�E�7�6Z<�Q	��݃C�ʮ}��@N���&@�S�J����p=Z��!�h4�jCV�';2��d�S��lp�� jI���1UH	�8i�����v��������{��e��;�fk�}En����n+#y���xj�Ʉ.���o���I7`n��N�+�5m,襖�-t�0�[rj�� �Q��?���tӛrm�5���;�n��N�߄[�׆���C��45�$V�,�G�˞�XK�s�
�6��xM;f�9�}�+���BC��.��-3k
��tY��,��h�ݦ�'H�s/8������r�IzlN�� �����R}�~����mo��>�G��|.%-)��h��@���od${%�%٣�d_;!Dq)*{��^�{���EVY%ܲ����+��{��y�����u����<��眷g��9�W3�����&�mM8�6�C��='�p,�(��JR�U.(q��x8FUZ�U�<[u�tz@��Я�b`(	�l R�M�J��ߏT�\pw��f����G�̅�-c�~�7-pݴ���ϧI"�tk�F6��0�0�î/�>�p�Ӊ)\����a/~l�f��~�*��ܝgu��78�.�w�/�T��<6���qtF^�n�m�>3u��O�*JVi�<2��<��:x*&O^�~�Emӓ\�W�a��mb��SA8U4jÆ�2\��7\����R���t�όc��L�ZFg�g?����zB�HK:2��Ԝ�e���s[m��������=���^+�k�S�ELq�����O"�e�T�Cd��~�X�����)a	?��N��d�\L�FD�=i]ۗ��"��{�H舨tP������EYK�4|⢶��R�ǀ/5f�ŝ��k�*�>�˯6��IJ�E�O��s�X��v���1ST�qi�����b����-9�9���FĄ���:����zG�lD(�g�1�&7�dbu��4+xT�����[���#�N�՛�g�z�>O�uHpݽIq�{Ӹ�j��t��2/�//1&�7��^�ī��ɧNN}������Ș���O.W�<�o�;��B��0��0��<M�74�GÑ�u�W�ߢ�W�ا���_����b튍?�437�&g@�._�Nq�Ն��l_�>f���).�}�Ƨ�����֨29�;��c��=.7=�E���u�n�i���cX����M��t�9r$f�����܈Uk��=X���c�8uǬ{oƼ�O'�}�)�c5��'<���%�z�����O��N�P���d~f���*�']VG��yg+56���2.3y�+�qwIH%0�m.vN�V\�_c
 �E���Kn��ؓnBO^U�٭`NVRGP��<HfE|YE!��?�̼��Eʿ��:�����G�}�ʂ����"�v���
$�f�k;��tL�Y�V��0|SU^��a��2n��m:��*6S��=�'(�>�/�9'��Eh���� "_K ���)�4@���g�fN������9c���:���3��w�U�X�*ܑ��*8�|�`�c���!�jzk[�ƹY�C+�$���8���Թ[58W_�1�=����|��,t������s�s��-�}T���ud01���VVٹΠbT��p0/-Z�	�7M��H�*GXC�=��㵩�!nW���&��v�z������V��fZV!�{��,(�*�o�9������*=Ln(A��e�yë��q�V���ue8q}�r]Kvd<���:dX�k���J��v�G���DbiMY�t��Ћs'�tz�AY>!a���C(�w~�����=�B��^y��9����܌K�Ԓ)�0�����T�*湟�2VӃ+C�H<�YYD��e{�>��Єp�� G&�����sl,m/V���ح�G#�TT@��QH�������S���H��5�tOqoa��'s7Ї�P��Y��B������������M�9%�b��kp$S�AH�V�L��@<�r�'*�>��	���J�~��?���,Å���q�B�.򓟼�Č�P��+̥�y��"��|�JuW�
�'��i�����:��3U/u��j��C�/?4�����uI���2y6A����߬�Fw����YzY6�ޯ=��� l�/3�gy��4�0tW�E�\�׿6��a��6�5tkI0�~3��с:ܤKB��*r����Zg���ٿ���R���X�������+Y[h$�Ҋ���	�NƔD��J�>����N��׿�~=w;�W�u�C�����
i��!_"��6�<+��.�������rS�?���G�4��Gާ�}4�.���31��Z#	�-e��@(	Ȱ�<�57�{�h��|���Fl,tf�Q�8�6��ݦL����y�,=��Y�3�}�2�:�N�ۮ��,����a#5]�d�
E�[�5�w��^���`7�N�c��9�˨�8�7y�}�,~���FKِ^V�v��黦���X�(v����硩��Oh���em�9���Q��N���%�r�����&�]�\��}q��~�_2��=�>晎K<��3���
��fڲ@P"��RiG)$�P�9ԥ�-�m��2�[>��-?W��@4oܰP������1����=%�8�"ب&.����������.��}�EG��_�<\��-s������L���
J{�M��ߺr3��R��/�Ix"u���Za�"H��<���vv��z�H�!������z����
+��)�V��V�SOD���7�җ3�Ru&�����B;X�=�.�~k4?� \20��X��Yf�Gl���P��
����6N`�)ծ�a9j�ч/��*Won�f��G�o�<��=��Gi3]>���M���W�X����zU�)��o��I��7�Q)9�����^�k����b�t�5"�������>{D��	keQ�3��z��Sr<�E�T-y�ڊ[f������J5��Vջ���e��H�V4:�gd�C�1&}mhc�BX�>�)�5���juDWha��Qˈ�iτy�U�<oV�=����2p�)��B���b ����a�9���m�:�	7�~>�H���� ~��x �a�E���Ϯ��u��x�򁅩�d���}h��%l{n%��K׎���ˆ-]��9׎M�f-9q���V/7Ewgc�����w��׻N7!�!��{e}���b�@�x�Q�zR��J�Pj���oZE�؍�U3xu+�7�a�J��fbuo�gD�*��9n�p*�;T��$k	������r����4ҝiu<4�.��-����:���Ѽ��RV,�k˯�sx�M���񅱏:<�����m�c� aN٧��S2������R�t�w�:Ad1��n�8��@��Y(��wB�fq'TE1Ou6��֪��H�H�~��X���J�M$�$'f~OEr�T]�As5r%���H��\���B�Ϡ��`��͙|*/��Ĺ����<U<0�B��W#i5�n��j����3( �j{�T ��~R3���e��!�!J�)t�)+S�h���v*1O�|�G.��Ă���٘*mr][C6�ׄ!j��x��@������<[h8��ڎ��)�cW��Jf����I��T;������XĴ�������,4T��ې���f��	�K�G�L��nF �-?!į��2�����<&Mb�ظ켥�V�܊�&��KVl���{�7�h����bL��{���&P���)�ރK-�Jn����Mq#��}�sG~vU�tO�~!g��~�%��[l^s�ǌjO7 _!b�+�ǅ�aC[���B|��q��M�ږ\����������x�7�y��o7��X�R��;&\׮��c�q%云�ه?�-d�Zή&�Gl����]���8eŖʮ���??��8=���gE�)�:cM�3���N�R�h���b�9g�V�j���}�(��=�M�|\����<-�8pg[3�B�GU�V�O
�`�2uK��/�̇k����B��ra/]����w�K^�q��N�4_s���G}��5�]�OL� 4�(�>����L)өz�x�ʻ�ew�^�+�i>�:6[,c�S�+�)O��i.�r�&�3}�49�&"���/,saI��}�>�����.j1��:AgWq�ءN��Ɇ���tԝ� E����6�)�p�F
��G+�
%���Y�7�c�,']�f��N���Q��.$y~v�|��$��u���-R�:ߟ�rS��W4�M��C@v�� ��Kj�tq��kKbo��7��S1�����\�]��μ��Y�=G����ɹ_\����L%�R���7�e$i���&���Q`}�=�ӱ�b�7ZbQ�Yn�wAr�<��!���_�7)�W�>�?	�ӎ���Q||+c��@�~q3�9X����?��5h+�~����6�{�������dX����ѧ�Y�[py�[��}9Ћ*`K�Tg���2����O�R(s]@(��s�sN�`u2�����j`����������]6DmOշ�6;툒+v<�a��?�S�p��%���u�@��}�0i#w��a���,�&yH�e��Ip)5snF��.?��X��z��W��j��EW☩�/S�����>�k�;_	V������B࿰�K+Wr����s-�.w���>k�(��#_����?w���MR�X�ֽ�H�3zw����*��#X�E��_�)-��ِ�Nb(�&/�`��ݠdUIk�58���Լ�l�A��C�����}y���/�əT0*!+�i�&1������i��
���W��vj�����K��n��e�Q���e���녛"���(�ԙ���r����\�X�'��u	�}��lx�Fni���K.�Pg�=��90p���ϛ3��JɔU���m����|���@��ھL������%��g�|h�V7�ș�����Q�G�좨˲�����n���{�q�
DB�<p�`�R��>��m��Bvr�{�ZP�f:���,r-�W�&�%�	0�M �ȏ#�
�xD����:��F��ȫ��E��\���82x�-�"�?wr�u�w~/�AE�[��mu�/z��Ş�S\^�j*�E��}��aw��=bo���z`5�i=���k����;���`�3���ga֕�/�|+��y�S����n� 9O܉�t�OGh�<qk1{�ϛQ�8t���!�q%G���TD-�S�[��!�����A�ŭQ���8@q����n�َ�����d����mb-���>��/�1���d��j�]�_����4��Sץ��N�ݴ��E��yY�����we�l-51���6;�]�1��pɥш���U�ŧ��rBU�޻������C�vR�e�U'��Z�"�,m!HVDY(KZ�F��(#�,��=�����!��e��=>��VG�����#O4�ׯ��	t�	^����S��[���J��l>DD�H0�s�D�7pM��u�����t}�4:1Ӵ"IˏR�!�OW���MT"[�=)�i���5i;�bv�U�J2����� 5�+���N����6��J�\�o�W�D��mF*t���0�w3�2��C�%��X�≎�U�Jg�����W��]4���m�1�b�N��h��j}<�#o�͊��8qs^��"��(�������FJ�ѦeR: +*�d�`aDܩ������>��؄��_��2܍�N��Ħpŋ�� 2��'����P�f�
�Tڻum�yyV�q����m{,�W�H��}~�H�2SknQ`5�b��Hr�]؂���?ݞ��^C
8`67�o�kS��k�%��^Dw۱Ci�a8��� L���f6%g��qX\�[���BJ�t�+o�K.F|�aV��-���=�eȅGs*�B&�Nq��i���������咅_�C�۲e�!l�
H)���f%yw hN&ll\����[$FdR�y��6W�g���,}����ef7"�U��/}��!�I�,����d�!�kn��РI�8�s��Ӯ�$��Μ��΅jX�������tE��y Ac�
��Z�	�@���e�E�R��&/�L=lks��5�>�a��&�g�<�9��+j��g�b��=`�#R��*E��y�T�r+(�m$�$��o�Ջ�}Y }I�,/��k�:̺V���JN��DxJ�ch���ר��Y����^�LJ{���2��0�v��{�'џ�2�f�M 	�J�&]��6��K	nUx�c����

��b�#���3i�Y\G-����4ܤ���E�+�:�p8�_/�16�LcKz-��_<d��b�Tn��*+Rs��uOq>�$F���O���'k�s�X��+!On-���5���`F В1-JL�Q�z_��U���M8G`5�O��%>J�\˨����g�Ze�x�~H���!��p�D�
����	�2�]�i���Ւ�p�f����C +L�4�z�ϕ��#���P���/_�xB��W�0o�������rX=���pϷ��x+p8P[���4ٵ���M56�N�����b�& v(2�<��uv-�|��k����¯�Q���e鄥�fK�d�F�d��b=��C��~����ձ�ψT5IUn�?�5Y藀n|^Լl���� N�*��D� <8F��q|B� �;G�GO��/���Y:�5�NܞUuՂ��#F�d�EY�����v*m�$w�=,��s\=54r�d7�<��n�5�J��$��$�D���,3�ݞW�B�Y_̿�� �m�b.���M���[Hu?��(��-%;N�
Gj��K�YڵM~��+׺�K���h��@"]�����ƽ��a�7'�|��vC�/+ą��b|��@?wWK��+bҍT\W�,���`�y>F��| u�@��O��_�����lX%!���6{��B��S���Ǹ#�u,�qX-V��i��j`ȿ\U�!�"1�̢�"1���d���}qd$o�ֽ�I6��t��~��kd��</춀�E���?������J4���o,n\�i�~���u�l�<n�E�˲���sp�#�0n�Q����Q��6Ho�����B�W4�Xn� ��"ټ)mF��X�x��֩�Q�nyA���绝�aP 
bI���/�U4Y��X��q�d��X�Y��\{y���c�y�>�`)JVtS����1 ��&W����S~W�p�:p�	Y��cF�'����i����X(Hm�Wܻ����^��k�n�v��o�Dς[��A��j\��B���'~�J��Ym�K�I4@il8��L_:��%jw��o�0T�~��v�d��:�}�]�2&��ߥ'�vn��:*;��O����<Q��hNݨ����%b�*�$9�c5L�`iz�!f����h>o-ia.�Zo���X��;��"�(�$�X��s9�׉�
"@�m�B�w�M(�� .�d1MZ|v��!�?�s��vӱ:���((Z��69?���<����_�j�ɳ��2�,0l��t1��n�m��EÀ0	�C`'���p��� �	_\�,�$��Ȏ�����6n2���b�>��w,�BÆ��F��: ���#�x����lMg��sf֞ Jѽc��G�n0�D�9��8x@&�rmH�D�N��t�K}~�ZI�
�����ѝ���'��YV�rI��*H�Ϳ"_�}@�aN}�U�hz�q�����r��������+0��^���!�u\��	)�Mcɧy=���✕�ָ��2��3�6 [8#�c�˓�R��lH��o%�5gy�V�������f�j�Ò�{���d�9ߧ��R��^�f�_�߸0V�5D���\��j8�$�ٹ�|����j:���pOH)TW:������+Ê����y9��񚨝��W�>i;�ݴ�~�k���F�C@CDf���r���VxC�Ȋ'�A{ۼ�p:������'���' ����P�5U�r�ƚ}��*��q�C���~�cp{a�E����&`!j(g��>.8f<��xa,C$���6
}Hk�8U�臨A/�"=�z`�}&��Ԇ���R�X��gǾh�a��b��jɕ9�4��>��R{k����b<�����J&*)/�O��?:�N�A��VsZ��c���+,�����;��zb�g��QAf�P���I��q�����I�����W�ІG q�<*����v���z�:>Nu~�@,��D�RذL�@�]��-��'�^ݺ��̽/N.�ne���E���c%]/P���[��,��1��Iƀ929�Ң 0�y�8�:`���l��*��W���@�h�����,k��z�%�<���x+ �`�!f�CI Z�r�2���;�� �!�0
�L�Pц�mߩb�TZe�މD���Z�@m	 ����
��7'N��=�#��9ߛ�g��W �k/eW���X�[F�*�0�7��ש"�zy��0>�{ڞ;ٻl��sM�*�A��p4�)aɣ�
�h^��G�*W�ٸ��_�Nm�Q�n�&�>S�D���_n��bn'����Lx֌g`V:^MS�.<�׵�o���v[q��|�ǥ�[��l!�L ����>f3�1Ε����j�=q�-m�b�e P�W����|FR�;Cgz	�u0�!Vz�,�<���6��I�x{�� $!�[|m]��J�RpFJ�RQ��FE�|�-���Q��5���?��v"i���D��P~S��Bl�u��
M�D�9^��e�<���I�Pp9��@�jDVd��D�F˟:B���'^� P�� ����ܞ<���7UMr[h�ST���c�~F����k$�=0EV�̾zs4��~���R092������N�x���J
bå�[�{>,1�vx5��� �����uȥ�������\!J������٘�f֎�_}�`��Aܤ2��2�K���!�x.�����⾓O���)P���Jn�oJ2}u<�a�Ȏ,�i��g��w�\wo
�-���<oj"�͚upQ�ټ�Z&`�����wR�G�6G�l��D�����'�v��Q��H2���fŏ/�M��P'���޺����t���/���^2�1F~��y��ku�KZ*�{&��g�"���|E��wFQTI��{����uA��ʓ{~�`�p`���WFD�؀�ڒ�^[�=Zt��D֚p����^�.����Z�D+����`��>}�]�IN�A\_TK�a�W<��+��ǗN����.W�3�R���b�m�B����j���&�� �	~��`H�܂p��>���B�&������de�}��|*���M4mt_gץ���+�Iwq��]�~����-6"b\7'�HA�<���C�tѤr�6[xO�ex��]J��I�&�t�n���_Y�6���B������d�g�F�~UH�H,Vٌ�,{~]c
��}n�4৐���a���qM �?�N�l��l���w��Jz춅g��x��q�4�{S)���j�&��;��miܑ�1k0􉒜6�}��.(�tX�������	�(+�+�tv�I���W���I��a�;��2�~�j��~q��@A��������ۓ������;17 ��|��q_����
��gG�.^=eE��􃅃���2jImq�Ӿ�Ž^ã�Atn������Ws0���W����DM��P�}s�(/���t�U����D��	��#����8f8�Ʋ���a���,��{�d��NTl�w����Q�����h��O���j����	����||�` ������{���tñ}ڠ���ND� f, �����q�x�ǹ�����&��z0����5u����a�k1�(��������]zSʓA\�.��&���w�n��G�"�1-�����%�%qIn�����I���/*�#�t��z�������<A�p�A
�H���&�4Hsڤs��.u@ N bs�X�����e��b�Q�	E8��T�������L? IS%�����O����!�<fW;��>�ۅZo��F�Y���Q��-���~"����^z��l]:��$���F�Oÿ�������&�@��i6��I�?�"0Jբ��K� R���rڇ-���Ƚ������aO���+��s"L!�/�g���=�����)t�z���pڻ�:L������'�9`	W��{����ꦔ�����l��(�⻛���������ݟ{�cQk	w��1�ࣕt���*�rG%G��|Ґa󇓏���ka����}��Yx ��4�Q=�T�ګ�u��C����[�� E���gKH$'�����>�.��7~,:��Q	�����n�d��'%8��?��c�c&�q���cF�j< G��j<��]�:�<i���q>#���,DLH+RG�d|o�ƥ~�t�����0���ߨ��;h]����|Ͳ��'�ȴgG^y� J~�u�pJ�2�֠9��}c�+;���L����( ��y�wD�\r���
Ե�f;�*�a��k���o��:�|ڮ�f1hp�C��~��E���mQ�sM����ɉ��R�R(�Z��x�qK���O��b�'|� �x8�����+��'�+�2�:V}���Ӟ���[�����i�5]�1'VEe�x09S%��^3<X��������c�:�wJ�97,Ia ���uV�Cc��?V2��A�KSs#2<����<��W�L����Tm3���o1Q{��><�r����V�"Ӄ�~VkqK�cx"uA�39c��	H���7&��m�/?�kt�1J0�@��Dų/f��ꏟ8������q�%⨚�^�����@X�q'��_쑍�'��L޵x�E���>�Ņ��NF��H�:Ę!k�7l�O�1*�ȒE�CI,gw�g�MaK�ڃ�dL�˃����1�����N/������?έԔ�P��C�Y��K/�5�L>�&����ҴwwB�o!��c��P��!�౑���K�s�l*�i��H���·�����*�Q�e�Y�[	|7֘Ұ޾��څ��Kc�����s&⓯d�E( u����|��e񼛠��Ó���5�-��ߌ�8��)V���,w�!A{ЖMM���*��׍�8���r�_��"�m�qv����u"#�� .���QN�a����~g���Ω�T�3b�}�u���bh����ue�ROM֯�v��O4�����_C��Go��Wp��OY|��_�	�5�,X��F� ��x��:��ե��;7�m9L����ί��Җ���t��Y�p�"���X�E8�)��_����qA�P�}~��N k�����Jd�忹)���j@��A����_%{[j���X{]�ZZ���	�]�=ok(��i�hõ��*,�Ȓ��n$4^�����F�U�|��&����7P���;�βw�]�((�f��i7�m���5�o���4'�ʽs{���y�1��ˡ7����ƥ'�=�d���=��	 ��'�q�A��)����c.�����b�����#�G���kC��XIf��/��M9 Ǫb�S꣯T�Ͼ�o`f��}�����yU{-�\�%ֳ�A���?~ �&1�S�\{�W�R`��l��>�z]�e�jiתݟ����d��5�}_sd�|��N�%jP������,���!Fۿ4z����؜o<�o*��C�7��R
�^n+p����y�	���P�ĩ;�)����v%S{0ئa�9���-4��k��-G:�
�F	,Y.���#��������/0�} 
�˝<����?^�p� ",�ةD`����m��Ll:�5�/�:�3ɽ�~������}�(1���ܕ�g���'X���Y�2c��	^��|���Q����Z#�w�(����Ol�����^���f}�(mN2���+��a�r���|���Q(��{C���JN����Y�߸��CzJ%mt�xg*|���R��I|Lz967�C����h�����7@���+��d ����(�c�Y��ۊ c�uE���U�r7&F2�d@��B^or���:��	0:�DE�M���m)sq�Q)�K߶m|���g�*��x�����_�(��m���T����E*LӃ�;���6j<��R���Ӫ�Ã.��VtmFp��� ���Q1��(����I#�����BW($�+�g1��z����I�Xz�#��Ư��gh�HV�K�A��7?�Is�M�j�v�?�4�g�!{�>f���p�qSCUp�[�B���/�S����<������2d����M����r����^ͱ�VF���= WD݌�!����Ѓm?�U��L�J�S
�����)�*-���\�t僑��r: E����y(����|y1�?�h�&�{� ���'l%O��DSf����$�����X��?���q�.
��@��f�*@u��H���KL@���[�T[�����
��HNL��D��]�u�Aw�R����%(r�������������g1Zs�]U����Ɋ�^-euS��=�]�"�Web��C���o�������U��9&�h�+b��5v����b�׭�~��s�Yz��:�Gʯ
��5��u��4J���:%�2E[R�(��Ģi"�NQ=�v��v�]�ʫ�[�,�M��Uu0/��+�'�u�~Q����������Nm��X���w�bM;���q'K���� ��F#U��:��C^3	�D�������e��-<�T\�#w�ϩR�0�y��7bh��*U�!�Y����Nء���~�p�����=�T�jT�I����}�	�z��vk�z&F�����i&pvt���9i�/��{JC�	AN��-��3�\筵�f�D<��t�����,�P6���C��x:��@�Gj�R��#B����`O]� kX0�����!_42��me�ǴZJ��Y�L!#|v9ط�T<���7�}��A��2N_�HR���L	��yډ���m<0i1Dy5lܶ�Ì�=gbdz�l��%�a���ʠ�kfe!q�����>���мOb��#��y�����n3���nRܝ�v�x{�i�����.g�ʤy��q�}Ϊh��:�uy[������3	��3�u�P����c��%�����3�ළ{܏$�&	k���$E�K�s�kߎw�ą�?�`��F5���ܠ�z�L26��A����y��ڎV��|O}�y��U��(�+��i���5��w���,$ݹ�1��#}�Z> "��̬D䰤Xh(���.
) �>mY�S�e_�'�	�9��?��["��^�9ebd�W��-�U ��JBR��RϪո�����H��n�կ�}���'��<m�����H���+�ɯ��k_�F�)�y�f[[J���Dp��z8k��&�ӮN�`1� �u��c�Z�(�� ,d��g$����3����d���� ����1p��m�+E�F��}b�cЙ�QŨˣ�e�� [�u��Mn��*��XV�D� ��H��P�3�W*����O�Ŗ��^f�Ǉ�Rn�֍v�z�ckU+G���A�b�kh�fw�������L�&j�Yɟ>r������[�,n�ǯ�H�L�Un��w���\y���������>g#ٍd 9����>� ����-ߛ�0d��L3r�yK��A[y֎X<_��z��4�����:���Cñ]�f���V�R��o��@Dɸ����Ne��m�'�)�������a���Q�E}�ʪa�h�D� Jb-�� b��c)j�`c�cV.rpK=�
y������6k�3�S��$�6Z�.�D��T6��ެN'�i����;��W����>�.�Xu�T���������gܠ�w�&��,ѭI��"��>9tū�~C�ͫ�yi.6�=���U��l�,c�M�dF���#\*?/c��9k޸��	�`M�a�⼑&�+��	�#D���k��u���E����u��-���Y��l��s��������Q�d�K��[�~�=P�+`c����s���N.Z⦪4��|�_��R�Y�V�v!�1w�HhN�$V��z�_������� 9%0w��c�aW`��Q�76����f���oY�LP��òo������)���8ְ�&r �Xheּ�'�х�Vוּ�_J���do$l��*�	���$�te%E�5� ��	4��#+��˝�x���?<:♽.{=L�>r����������%WSM�)��]���;���V�b�y.`"���b4��="}'JcS��7��*1�S��f⨨'�P@ޣ��ŞaN����[Z��2��k���i6��Xys���!����_��:��ٮ�>���$�X��-�1an��(ٟ٘�G@c�?_���<��o�w���Yà�H�p+	��m�G��zl _�{��}�=�jNj���z��'<�*4�����3�1�ԔEՁ�E��Ҹ�ՏR=�%�����?]��;\�x��/��^P=�:Rs����ԅ~^�tio�*��(o_'42Ɛ��1\�����$�-ɦ���l,`*]��O�6��	�V P�����������uo�+�u�\H&�	4> D��??-�8��� �e�%���I	�s �[v6z��tV�Erq�/�����FS�"ݽ$ �{oO�^ԑ����� ��w �V\�q�}O�u�t!_��4ŭ�.�x8B���x��R�å���A��U~%��N��Ǽ�������;��"�g6x���2q���==��4�@�#F�7�/�Z�D23?>�9���߃�6�o]KC�^��[���O�X��k�7P\P*��@�NC|ڝ!J�j��QGŏ�
 f�چ���ĬS0�bш(�\�c���&4���3e��ί�R�r �[�Zע�jI H��%e./���y98�i�qQ��S��%��TX:t�1^)j)4�k]���G�"Q*�����D�����[<��T�E��й����DזB��&��)�܃���_��T�P��F��ʃ�p��D=�1=��=_�0�T���ܿ��̋W*��������&�C?�t�.�n�3|5݂W?���7"�rs}䇶���d�!������'@������MZ�<�����'�fTQ#��v��Ύɵ�Pۃ�/�\X�M�~�I�)�'Po�ku� �,�;gI{��b����sH�au5I��M��E#X������\�4��GY<�IY�ju�l�y�$��� )����쯮��x�D����qN��F/EJT���v�]�p�+PB�#����j-��M\_P���|\dO��y�
ȸyj�!�����;Xt���W3k�1��D����*7}��M�<w\��B��3s��ub�?�����$稗��񺱴���:I|;ūon��	�?�iV���
������E����P��xѸ"�yp�:_3I�v�u]�bL�A�n�j�+t�ԷjH��������/$�1�o�*p��\�����#�}�0��n+#��+x�8޳��4�2�0��@s�E�Un�n'��4���7�q����S.�N�0�TLȌ[��(�e�%]���+�#����z ;��i�I��x�'��)MJ7��n3���4��|o��Z�J��4D��^�n��݌��	/Sj���\��'��#�I����u9Z���L�B�es�����?�e�����p��1ە��O"KU0`�^6bF�����`��n<IS��؅k��6M�ka���?�g����(c��A<�-��z�@�Ձ��e�$ʞ��wVEH�w���/.����o`�"p��� Z�$p<y��7�-/u�P��-@�T�=v�_M�vU�2h��귡-+]~�@��i�y�9Tp����SEx�������z�{�@��_��V�F3LX0��s�Jp��<d�]l�
�����F�9��#�./>��HB;�\Z�ؗ���?�NߟI���5��3�A2T:��������Jz9���^V,t9�ܥ.�{#�C��i�p�7�+_��ux�N��# ��*R�)z[r;TF�@;(����'��p( ��zM�@wǨU�4�B����ϰ���`?n�����Q�	z�.RV�捡�7�g���k1�zm�/6�T��.�=�ϫ�Q�� ����?7t{���[ �u/���꺴���	N�m�����7h�K���`g�|Va7��y����ítsy�y�L+>{Ի��͊N`�������8P5Z!��c^Z�Y������C�t9�rR�^��Q�ok1d�e&��!vC��C�m��Y3�_���O��~fg���,[
w�����Զ4 ��x-�H������	�A���U� �t������y�O$�Q���!���8}���W��ˑ����Y.�dk�&&Z�S�S���T| ���x.���ǋ������c�d2�HD�xQ״��t���c���o�v� ��^�ʢ���
�`R{�Բ���L�L�#��!�}�����ʚ���X2pG�Y{^���B�P��i�׊R�'��	��70����x�j�ҒJk%hC���vU�x7���qyѷ�n��xx�aG���N�*oJ]'��E�&'��~	��p����W͒΁S���Z��:z���6����j�\.�4�18�^��@`&DH/����%X"$ � L#�$lίD�@
4Ps��oi�WT�Y����+�a֥<�pRk�6mdլ73-"��s�J�D ���w1���ee���}��b~*�*~��1�1�W�i��j��>+�"�����j��Q��W,�9���-�P�Q�ZwūH{Vb6~)�����}Uę�j(��~�*��gO�'<V��c~�d�~*:y�7J��y8��&�0�c
�,�[��w ���f�]�[���dA�m��� ]U��W��Wc�cV2�QP��y8gA�w~�6+��E)�����u��3�O��rO�+�
$B7"��|�ECl�$���2�'���q����C~Ĝ�C�姿㘅��t)���k�ޯ=��f�j�G�ᗼҎ�E����εH�����^gy����3�^���`u���>����S�/�$l��įX��e��z��'Y��Q�=�I9��o��z!��ָ8R�����3��yE�I/'�c���?rlr!�p� ���Y��h�,t����%ɞ�����Ȇ}KwC�q�>Z���낼��et3}V��`<v�lۻ	��(4����	�!W��c�-���SaY��������}V�zg,D�&��� +����Sh�O:��R��y5jP�x����B+wr�||>�J�\� �3W�l�k�+I�\�*����V��öJ׈����kT0��s��_`�U�_���i^`�>��z%D��C��5����6֝о�oL-����'.e���A"`����s_(����n���5F�W:Jq��g-�v�������U�m��@Q).s��7����k��́D���)�44�/�V���Q�EU�r����yR�-�.-��d�o�7W#�;��X�ނ}s�|�ʈ�`��m[��18:e��v�7n����O-�X�ۄ�m �ۀ(s����x{�	�Rp���6;������c������BZ�$JB�U�}�6�dg����D�����#�{d�({�>�c~��}����~^�H3s]�|��rι�'9:�{�,��2H� �jr$h�i�"�Rd���!D����E�i��Uמ@�ƒ�7�,�u�W�'d-�����Uz�^�^��Vh�����lj�v�ݮA�!r9�z�m�_I�t΅��A8Ѻ��>Z������
�?}��4��:�����l�3����{��zLON^>���˸�R��wp=<̣{�l���S��l�{Vps�F�$����l=X�N�%���q��=m�1�9������.���Rb�����(U����ӳu�>f��?=9|�u����ؽƘ�E�vԹc�z��Vl��f��E�����=1�ʾ;~��̇;�+�f�lA�5�+ح�/�:�{}�eآgȤڴ��v��`����A�j1�3��Fo��>��).zkqM�q���={���S��R�:�O'�5����j����y�>n�B�=Ѿ�]z�Y�������c�rIjX;�B�f�Ng�/M�
�-�	;�d\����OpcQ��O	��y��Ȓ�%N4:�?j0x��W�+�Wm�~ZcUժ�R�'Z�u�D�5�wn8��l���V߅�
�4h�A���
	�����U�/��t�	������	�AHN�bś ��������8������ԝ�-�h�M�#�<�UWH���'�ӵ�wy1B��0��g�&'�����jS�"�K�9ʯׂ�K�hK_: +g��n{4�#��JoEލwj��:4�E�1?Gy���SIu&^��b�b)�>��j^Ƅ����;��X��1fY ���̵�d��ӹpF?�ֶr��]�M����d�M���(щ��; R��,]����V7�+�]L{�̒��D;�Q��9��a�e$Zd�n�*��[�G٠��*��-�𫞾�jt�>��*0��9�=��>�{�`XF!�o� �����9%��s��J���"�4ц��e�%��5���=�^M������P���D�v�nE�=�`��݀9Z��{VS��'Te�,n�H����Ҩ��W5��L�6���N�пe�a�]{v����C�M���}�0	9�����y��T�mCW��#Ϗ�M-�t'�:޴���ܟ���ڟ�>�h#�}L��M��~?�T��۽~rX`����
m1ɳ�?��c�b]T4I�.Ly�p�1[x��H�o��b����s�fZ����S�c�B�D�O���f��z�m[����$�a#ha~3��Wa����o���1Tx�-m���X�{��]�����8�ٞTUONoǅ��磎䳯a�d\�����ʕ�I[��z�K6"�qu�XTjQ�r��R��sR3rÝ�����Gv��0�j�x:5��7�#���e�;T��4h�]W4���ɮNuK��_�W�q3�#����U����Ō>�6 ښ}(dYb��a�ضj�L�-�*mr<�u�:p3�7�B�m���{ c�R�5�����V�J:L�0&ᇳ��U��f���$�A���q&>�?6�"[�$�?�l%Ulfx���S������mʚ/4[����@f���n
SVuް��v�}H�k��G5�0���ld�z�=(	����y{��CB�<���@���I�/�ѕ�W��WR���*7\�^���3�z�|��յ��F���?��o#���0�';����%�����$�5��b�r��<?Z���e��_�Jk�zs������d6#r�/��&�7�q��%,|o�u��>��Y���d H�-��kUV��*"�������������\�3�}6[�3������b���G�%�s�a����-���0>�yY4�¸�ɘ�ج�H!��)%�sG��ʸ h�o����<����{��Լ�ú8��n�!(o�](i+0�S&Z���ʥ��v<H��1��I}��|���V�abW��{�l���O���cb�_>�J���\�T��B�� ��Y��iya���Z�E�F{�{ϼw[Ya`=�����3�?��.*ⱽAI �/��Ϛ���ӖM�����d8(O�z��B+*'��4M��ƒ����~Ns����`������H���/�<{q{S�FQ�W7��ǚ��6F�����]��U@?�ڵbw%y�#H)T�SS�u'�{yZ���뎋^���|����o\�f҃Z�m;�,-��>:�ͧ�����5����G���"D�gv�hTl�f�`rm��S~6c(,�-��g,,�]y�G9|� �#��IjZ��o�ƈ?����X� )�{���"��S�f�a�'r��O\���7��qHd?L-�J7I60J�x�8�z��[�5�V�靅*��_[K�u��.i{�c��Y��@�~�y*����Xg]`ޙ �k�m�1������V��>���r���1����?��ڳ�o]����L�IJ�����E��{"a��<t�|�����*}Ђ�W�һ		G��i������x��'����9,�E\&�>�hf�u,� Ys��a�Q�R[$���W�M,�*,kS��}�x���BD�-�}av��F�i��|Y�~��j�����[�GÖ
q]��&��C�d0J�I���E19�F����ϲ.�Z�`�?pOt�qԘ�eXt�8]&����/[�5�5�S�ǈ��**�^�B���M��--�����ѵ�K�nST"�fy���U�8;�/�LVz� �C|e�P?�EM��Ox�!�|��������5��1�Yz2}�J�:��"�ǲ{�0��_�)e������<�GL,%Ni�O]���n(X̛�5~�Bg���P��Vi���n
%쎹׸�oѻ�~#�N{={�	k~|��&� �QB� 3��pt}���~�
��CP�0����Z�%�%A�Ř�Ǡ��H�-_�X~��`K)�٢XaQ����yE:D��8��awSڱ�m؃a����tқ�8�-��2= �����p�#���Uf^2��1�b#��KU
V�ul�B#��_.m�&2��}�jsM��h���?z��<������i�,��jn�{v��;����Е��}�e4���%��鋎^5��ΐ���9�|-�2mvy������U�GlO��~����8n�����+IT$�~K�y��:m}�6�(�h����MF4�'����kU�?4�V��2�sz����\��2"�i��e��wq�|�WqƖ�FS5� �0�i�t,���'�uk3A��xB�����9;��p���5I�C��Z���~����n�����G��6j�u����|p4�"@�\&!u���S	Jط�
sƉ6����U��]��N��:����~�͓r�,+�+�N���!=�����)C�g,���}�U�������+>e��:�Ļ�-J�����fZ}k#�iC5�D���a���ٻ"q��عS7�r��a�&>������m�����K�51��x5�?C�; ��>w�-"�q0p�/�ҝE!��y���+,\l��>��(b؃G��w�x�l���)/cF�u��Q����l:���Y|{�� ��* �3��a��+sk��;��+1��!Ů��bR�*��,@�x�{�Yd�7H����Ö�?��b�1d��kr�u��`3x��`�*����ط���1U�,,�.xU��hk��<{�fա���z�j�{��˂�*�t@l��&��58��e�xс"*���� *Q8�&�-'�;��Aw�P�,T%�P�g= K��ۛv��m|2Zo��"���W}��d��Q�\ZطԤ�3W�=*򍫕���>m�����"���-���= ?.��ۋ���-�i�]�b9n*��U��ۍ\Z�)Rp��M ��?�M��=�+�si��vi�\e���U�f���-�ei�C�
��
�U�s;�e)'�į3C�������{8�sQ�I�~�J��FK��������H�,^�� �����w�ޣ*� �7�.a��h�Gz���@-0��� �#�fl@z>Y�.+�D�1�w#_ڿ�� f�_P�;�i�����'Ą�Г���ٻ
����r]��(�`�A�#����Tni�{�Oa|K������O��<�֏��F3�V�a��$
䛖*���o��.���j/&vV���D;�����)&�����iLB��
�R�h"���>\|A0���yg(a4l�m-d1��>����ـo��A]{vqh�luL�kk/�/�q��J�Wdᠬϓ.����e"�4���")D��u�c-��ҳ�5X�)�!6���ӿ���y��I�q�y{p���\W�R���̀~�<Ŭ��S�P#���"�g�P��К���9)��Ɲ[�W�aNDfe�\�V(���Ix8�I�Hy�fF�.b,ùkm���Mjk����Q�'���y�jxv]�B?{����H�I���d�|�>�b��x������8�W\W�FZNk�4�Q���ԋ�UKO}U�i���j�B�P��n�<O��:�<���}'}��>ỮM(q�)��L���� �&�r�����F���J��;�.y����G�d����[ZNԌ��}���DW+�]%lQR�TKҐSgl^c#�߷,���<x� ȋC�n�����01�����.�PUi�X�T,��D��h��oY5?��<���QW���ze|ճ������z�τ�Po��)�n�Ӱ�IwO���y�S�C��S���UU��;YW����S���ޝ3g�JyV}4����#�ݸ�_=��C�j�o�2�,HvT�tq�ԇ����_�=��Z\3�lf
*x��N$��!���z�����̭��h!`��6����>�g�#�V�_�?*�Tz�)�������Rx�T����u��5���a?2�3�X����j	'#L�a�̔CǢH���&���lȪt���Q	û���|3�#�
�ي}��k�E���J^Y��ϵ������e��Q������G	˘�`�w}*b�����E�5��#qF��9�ha	#�=���K������\t����{~/	c��̌C`Ś�6���~||����+v�k��TƁՇ� сY��|wRh��6̤�ՙ<���)�y/(�^�l:��NR���t6/t��Btvh��8�{�m5���|�O�}���-�}�a��b�� �N�X^�����g�̄R^�>ޱ��;k�Ca�!\>�$"9���G��a.�۲�mi����N�X�&;���{�~�O\�ۚ�T��'��6���<Ŗ�~}s�{�8��6�!m�aЕ F��Ena�݃ꢥ&]=�Z�ڑs��mC��'6ʷ>K����o4#�����3+�q��R����ŀn�{�v�'�T�ځ̜8���\s�����	˟��A�x�N�I��+�'J�ƭUoN�$�&/�c�|��.��u�M96��w��� �Y�2��ɲQK�.�W����m��c���뽳�+�h�:/6�.�X/�������YEf�f� �X����Կ��gꖚT-ް�߻�p�ٺ�Җ��1XI����$|S弹WZޒ�
��m֑R�Q3À;a�.#���g,	[���?�x��_�-���8� ?t�A� �����*[�뽵e	�p1��Kj@?��ϴ�2Zu��#�������<�5L9�JDN�u���F��Ŝ)�\`���-"�K���o�-���d�FUf�o%�ǫ%@���e����Kƕ�Nx���ff��+L-��N(�b�l��c#�,h�����'��O�e��ri}[/x�r�sׯ���5Dטtꔹ/�&
V�>��1�����[�R�$�EXP7$-��%GQ��S�o�F�oH��>���\*��M|�u�w����(7Izv��W���?֬'S}Λߌd�RRD�L�n����OR|�(���������=��8♟^���Ͼ�]�TK�G�I� �j��Wm]�)���^	%���5���,�4l�� pw�=�B�=Ѕ��1��h���3�|��V%/X��d����T�J�W��e*|17a=�s�5wB�������4�*�lل=&��U������T�.h�F:8߅��f)��O?��5iL�4�=u�{����nۼ�0��� @8W�U�>��I�"7�َ��FQ�G_���mP�
����v�mVO����)��,��$}5�W��lH~w�v&�_�u3��鱗��/��d�xi�7�&1�O�N�G��b͏C�K�?a�kyC�tk�� �aK�
o9Y�5�>cKZ�8�Izh���&��#:�CgZ6Y2K;��q͹������a�P龛?/p��h�E:�L�����<��]��ԙ����+R�j���z��]\��]P��j����jޑu2)�@�>0Z�RA`BR���MR-e,}���A;n��_>S'6�`/�r>��SF�w�K�Rb�<ơ��O���y\q��u@x�ib`�M�W�pe���������q��y`" \���)��9�����z���s��I2�G�{��4@��/�O�]�@~�R_u$7_v���/��S��DƵ�=�<��� [�t���6��&MUy��,3�lc��x�(�mÌ˰򨙾�Y�K���u�;I^۶���yv��egj	����,�n����G�9�_��C�t�E��+b&q6�H� y\����������A}�Z��ʽ�C�7�y!�����N ���Ͳ���(�c<˙}���7B��'=	ҥ��lh�Tv��╗Ͽ��7�[�/�je ����B�\�F�53���F��)U3lzbb��'v)9�����E�0�)$�S�d�X!t�?�F��NE�����>�c�H������6}ӕb弬�@$i��~���^�-��Jj���?L��1�����ͧP��ttB5A�FEI�D�p�eנZw�ՂJ.����p6��= dG'���8x�찶���E�v��^|EGgac�@��[���hZ��(I���gs��� �0�ʒ������M�Uehl�#*���| 6�ce�w�%tތ����-y�={"^ؙ��������
B=�6�p���TK�u�*���$�)c\_�������_^��bf��|<��y��o��Te^�I����#���Y+�� �����!���&�cdT59��ް�"f^R�U�4�u�.6�h+��T����a��M�vt;��l�#`��m&��<�ۿ\�t�����Ja%��YX(�v��T G@�5P����J�S���q ��~h��4-��
���+ �pז�)AW��ޞ{�X��4������r���d��ɑx1zخ;	�������lVo�xHo^��(���9-y�	��Kj���������ו�cy��\k���{�\f[+[�F�S�(r��	�l��S/L}�G�a�IԺ�T���s(VVv��� ��&��ܲ���I��鵔�b����%r���0�F�f��Z��)���x�ɰ]�|�x�'ã���ٖ
m���8s����6��g쮔��
u���c�ѴW�!�ˎV�N��>�IYf
�k����ia�������Q���Q0��L����O����8���^K�W���jł)Φ��p�㔝���L��Z��]�M��F���	g���f����=�����א��. ���bY�h��T��2��{qA_:��>��jH����!d��X�Lֽ���#��ǀ��#/����l]z[U��=�΢��4{�O�$j���̈pv����5A��|%�L�NE���j���J��l^T\y*�E��/��{�(���	[Y�/�y��v�z��^"��>��/���R��*
i�o*2hl�������R����hE�9K�1���/;��Isz��n:B�趬��=������HW5M{x���5r[b�xq�E=�����U����U�f��aʵ��¢� +��?]�
�uf��ԡW_7��b?��";XaA����
�*X�Xr`I��V\<���(P0çA���<�=�(ɃG���@��I�0�'u�Ӯ�5A���ދu�kV�\��e��}N��`��#��RH��*��K	�$��_ђ�Ȫ��9�X�%9��[z?�Q�=F;MV��i�v|�Ś�1y(Ue���4��8yi@�׮�%3��Q��x�+p��I��@m/ X(7�xΓ,t_&�E��-(F'�r��z<�&���w�����`csl
�kp��>.�����\Zc;k��܌g벜2�C�E� aZe07��&ݒ�m��)@�<�Q������ZY��s��ԡ1{	J9�i<yR�����,:�gO�������:%߱�))���W�s�q9X����>v����hޘ$��c,r�;4>�����#�W��<���I+�z�
l�_ww~*��p7�R�R�J��.HpE5��o$l�K�d/$Pe"}����2T��� x��^�=�.t�>X`�n�E`x�к?H��}�x�ռu�͍tЇ���
Y�Dh�f�>^���n�WP4�ҭ��)܋�V���t6� �3�'�q�0��k:j�y��^�X)���yoUd �j�~S���b9}�c�#��|��Ŕ����8H%���H�m�;\�DXn�f+�v�'�ک�v7�B���	�@���43���J<ݪ���j�����*p�'���V
7n�>!��C����^�i7�����y�f���bݞ�qG�r�Ph��+]��ͬ��"����L���q!�]DGVl�k4�+{�W=��G1䚒u�zڳ��!�@B�K-J�O_���D�:���%��+,��u��_�=9���D�2?4C�Mw�	;P�W���j�&k�T���� �Ah�oύpt��̵pB�kn�?)���@^%ށ���B҉!p�}��օ���1��~8ڸ�IhC�3�]?|���w�O�aC��C	k� �*uZ���8T���(�NK��+>|C@����Ơ�bfU	�\�<.V�+�XD���8������XR/C�޽�	�0!�c1c��8O�DT�/S�	���Az4�t���.��u|1�����:�3G����o-RA
6�P�3D��Ą�3.� �`�la+�"�^-�
P�͠5M�S�[@��*��n�hl��V�>�qY�,��ڗ�^��[Hl�� �2ǏR(�;ק�o�o��wt�K�?�_o�Ϝn���r��CU�A����v�/�Gݒ�:�R���̸��W9�� p$/��װ�������nƵs����(�h��e��2��}v`}�i��g�0�Bnt�nix��74 �[Yy��$����5��(AM��+ܪ��a������$<�+k��l)	S$zg�۞1��*a!@���Z��;ǛY�k���s�Jƴ}�]yn�ݩ55���:��Ӡn[��$���$hk�(UH��!���5q���R��c6mUu�ĹD~���e�r0'�H��gV�����w�e1���2-"^<ގw�[K齩���oR9��*i��w��������aȬ�:�A(���7��C����7v��ܤz^�$<*�7��j��؃7t���m�^�2�3^��J�\��kޭX�7L��zd=t�+���! ]TA7D#p��v��Z��v�����X�YJQ��'(ɷ��ZRu�KMD�Ò��ך!LDʷ%h�x�=��!ݨЏM��<~$�#�S=��Ѣ?��b�H�c��Auq>�n�]J�������)��(�2�֓3@"v��ZWv0Ք����~CW�AV����|iJ����֞�@'c ���MժlL`��O/(�|l֜��0��;��!8�aIP�߽x�_O�Ǘwdǧ�P3��~�P�A:��=d�	�ѼTYÆ�B�`�n��9|�hi DMu�y��[��Nƴ�B�GV;�N�r@(t��3�v+��Y_'ag��t���6L:(Qa��kx�f�{��>��k���;�>���nX8��o���ǩ�,(4�P�!��t&\�������GP�]@�Q������@_��h�@G��>���y;��_;���j>Z��a0�]t�L�@�%3����#y�]y|<`�-D�[F�iٱ��G 
1Sk@��^����+u�������ڽ�0��T1sz]#��%a�,u����J�m�s	��7��2�jI[JP���»�XK�n佛�J+��#��k��Ō�����ϳ�g���P���g���x_VqEtƵf`.q���#�f����>n99xO�+�� _�(�S&��6Ak���FOt���� ?R.~tѣ��OO�y�M:�Α�(�4��<��j����>s��}�Z�\̌>�����f�*ڧM�	�e���d�b|���I�|�Zmn�+\]�ϱ� B#g{n�nsL�~#��O1��� .�T����a 2�J����\~�'�2l�u�ެ���n�Pqp�os`��^w@���n��;��O�ƾk��T��NmA���b��Me��b�i%��<�#^�� ��/� ���ξ�/2	�7'Y�}�i���Z���z�h�n���3&|�9�eM��E ��/W%ȁ�oj��N�}���y+�F��,�eAg���z��ڠԀ�X�_�aFV��{%/6 ��#����>�	�cc�˽C�� �L���V�?��w.������q����$&�|x�/7�����B�?����|m��}�3�	,�"�.����iH�_���Sbu�h�M�*X�\��Rg_}|��B-@G�Cq4�0F���Lq���_i��w�V�N�KV��Br��������#}}�G�)��<C�v���x�_ݟ�p|`�yzt�m�s1Q{�a�o[��A�����~,r��W)v�_�Y��(���� �2�rLX�+"hG���p�� ��^�u�.�Su����������J	����}�<x��y�GU+���0� Sis�v����]H�x.�>���p�!tw�Z >�+�cȹh_�#��E�\���Y����4�������M+�*V���?�����x��y�����d��E�y���8:kP�%����GkC�դgW��QK���]��N)]�����c�M�b.�)���'�ȶԲۛ����CҞ�2{	�3�����u�� �z����4��b�K8"������eC����W�^Ƒ@!8zF���>�h@���!�?�r�K9Ƥ��'����"-`�L�����M��tf)���&�`�k�$��ߋ�� �ԭ8KC�X�v;�!�LV~�X*lYЕ��	Х�G���'�<8H�#���=�E")�!q$�l~��' � ��qln�Ci�� 5�%y�v���C���R|�&�N�r�2�pV�aB@Tgv ��;��9ހƹ��ᄌ2w��$s��w�/�'�z�ȓ����ċ������a�i�GQ)��G�?$]����OJ�$��1�6��Y1�h����s���@`:���Y�}0ω���w�\�����Nm���T���2�*��[��@��(z�Tv�/=hY�
�)*' � �oA��)���u�k�� v8�̀�m�����V�(�{�]�?	��j"�}g*��T�S'�����]d䢤vTJM.�dh���O>�;R�fo�U���	��QaEP��#\tg_&�Y {����hp��EH5�@ B������P����p��u��۩t�o���'( �%�'�k��:����e3��8�me��l0��~̣'�(�`ܿ��WB�/V�Q�,9S �N��X�����n�u�1��Z�>v����_��0�K�?�Q�s�6�Pо���z3���KEu�A3�/����[t?#E��3�qe˂H-Mh��R R�gP<s�� ���k����vR$��ez�댼�F�:|�Ղ>�7X&B':�Y�	�ּŇ�V���ݛ�9$Ox^�"��w�-��V�u:��v�tm۸:��^}����~�e�!w4k���<]H.���1'�bi�N��1t(�h�	�?�}F{�S��I�.�W�M�����Ĝ�X��PT����@$c}�s�h�����З �y��h̽����-imp1��*��Y)�+���	�8�P�O&EAg�l���D\F��q����J�@�^��W���w�� z�{q��Ϥ0h� ��DN����d�-h�^+�Bݡ><���(���Ox���$i~�Z��t֒�8���TJl�)��U���[�wtp8O�M "
<?.Z/�o�\8a4J�xh�N�l�1tNO=|����=�AfƋ��?85T��t��k뢢	���A����o �)N�f�VE�s]s��+�/� e�k���_q��?�XC��S����+HvA���x�Z����#��9���'�|�V���Lg�5V�a��g!Z?֩g\ƌHė@3���A8�Hy�&Y���uҙ)$n� �@� ~���S�s���Z��GNg����5XML�m1��\��D��A�� �܃G���;m����f�[�Y~4xiK}���M4�8���T;��x�S��$7*���{'e�TW���6���@l�Dn,���4��"������qg=���X���Ai$�R�g!�2g�(��9 ��5q��!��G!�B��E�+) ��]3�xw�q��l�l<+_h-�X�]M֤p��A`��c�����4斢k|��S��5>�`'�rA���ߎ)癫�������s�-��	G��[S�$5�c�&�H�6W��D���l&���v"7�:�x���'�p�m�v}�!(1_�� 4�,贍ZN�"���Wi<Y����'NS�}�AE"�����9��v�pBs8�P�A�2 0-o�UGeȍ�S��q��a	�p[��Fk\@s��fµ�?���
�Y�A������=�t���ڥŴl�@l_�[�s��WAA�%� �<+��4��:�x ��I�l�:нв�r��^QX""_�I�dJX�l��AGH�����k�G���{��t�	�ϝ������n�����d"0{)���N���9W��:Y��Oy�������bƵ�6����O]��=9�v����7��k?_�3�y�1�2v�j:5&'a|'�@�Ż���@]֯�Ё�*�m�A����) 8�����+�v4/�gD5�;j���3�p�qT0`����X�����X��g��?ʹ�/�+��6��[w\���wW��w��V����G?ܮӅ��� �tA�+�X�?�������v.�����>�P�M���n�j
�`����U��y���-&���]�NN��g)���y�.eQ�Cg@��m������ADV�bkR�c���_��c�sIs�#��`Tд���yދ>�+��0�Y�fJ8�E�j+5VsU䪆�#�����q��,G;F�Ѵ��:/�*�Ѷ����T��tnAf]uS�If­���5������=�� �&�! ��^~����m���.8��~<�"��0u���	��e`�������l���.@����҉Q{�%�5gd�3߶.�g!!w6?�俈�:Nn�;�A;���p�m���Fd~q@�.0�8�r���V���,Rx0hy��@i~so������_�v�ȳC ��{G]�Q�2��B��~`�ϑP9H�VT�J���myz��GZo�e��S������ ��ִ�M�!�>�'# �H��;T�� ��mVt������YL(�j�mD-�x��Ś-h�`YC�	���'~��Ȧ�F C�~��1�@UVvdŒجA\�g��c����W#� �88H���˅�YL�m	���i%=�u0�e>y�]*�
�rz�[����`H`�nܰ�{9 ��j1�8���GHM�쇳=�)/ѳ� h9R6���N�O�M:}�����t���G)8.�9��M`�F��J&-]���+ͼp��[��	w��&����[@����;Z�T��~�̯���֑��C]6�.]��A���X%-!�J��6B��ol��rx����DF-�+� 4!�FS�oV0�tJ*4X����,L�3���r����/]���Q{Qm�X�9H/�¥m���,/��O��l�R�>���Gַ
�����:�G!��0�{��K�����`Ҩ�u0, �+k�b:5�����%4�Ə.V@����o��8]ޙ�6�W��=;Ƅ���V]=��X�����#%2�*�[h�����ȴ�&	v�	�S�~q MI��Tr���kÃS/k@�����R@�r�E�Z��IwM}5�D��t�j��@Q1��9�Mag�o�Cѧ5�9���������)�r���������v?fl�F���m�-�ϧ]:�Yl%8o���X��l]���~�B���M��0t\j���ӉR�.�"��0c)���-���QK';��<��@�����>���Q��T'���+qs��Jc@�\�W7Ք��_���uB��HC7L_M��ip�|E����$����17�v��p�9؈[9�G%����k=*������t�����d�l�j�~�`,p�?��塭�2\�����/����tN4�b�����a���̳o��m�����x��(Ӿ�[��))V �)S[�d��a��?F�����`4ARÖ��cz���N ��w�V�
>�8����ᣒ�3�@���n3�rvhu��!�D�2l+��X}N6�����U�U��cg} �F����E#
����ɠU_����Uխ�@)�Bo,,+Q�����.ݮ�a�݁�c�c$H���#nP
 ���H��[��tP���i���N���f�9��c�<G���hGJ�-C��4�} 1+�"4��UE ��+�1�|"��&i�����^5�>�M�>3?�}�\�uh{���O�|Ed��+%ԙ)O���/_���T�l3�>�v�U���Yy@�^aj]���r��A}�)��@���/k�~���|C��{J��Ȅ����$����6�{lAF�3"WC��fάЍ�������&į�tW,$>C |����2�����[�ڀP/9�Y`��{b`P��z�0�E9� �=%0bK���l�㌐�� u�U�5?�^	��y�Һl�h��d��-��W������L�=����|"��`�3EVl�a�"�F{w'�|?��Ϗ��>�� �ҞKL���&ʂ=,�6�M��W IȮ����5^UH��ސw
�E��`]��>�`{�R�`��j���b�kC���%PH�Wp�v���� V,��_qM�B1�����t�w(��w� �Pd��X��r���x�f���p5���sԕ�X�"��2���9I�l�É*����W24t��e	@C��[�Ya%JUf�a4�qY_(iM-X�sg7���H����2E8�%�������ɲ�'�Q5�����*�@����P���p`�1�f8��w�8ɿ[��(k��k��u�K��S���DM;FМ��ϡ�V���\��;2�0χ�/�Wb��y��#�N��
m2��9�K¹_��T`}�V5��|��K��ҁ�[�szK������]im���;��b�93�o���z�uh~�������vח;j�G�'��T������׹��4�++���?�9�J��x o�m�<�����f,�p��6�¹��DT;�"q�ܹ��c�.�\"�~I<C�uo/�!O��Q��̘Y=<5���8y��?I�+�I/D.u.��DG���^+j:s�}ؐ2i�*Ș��5˞�q�FŞ�("�ۧ�b��:����de��w����I��ڊe1z�qPY��\ײ���ΏH���pBA��#Z.���G=Ey�*b��|��ĩso���q9�`p�~������`��<戒[!���ν��y{���p�a.V����`�X�>x���B��Dghi�t�X�g�w>��}�#�˨cL���|�����dK!7�����Dׯ�|�e�6�B��"&�>_�!��1�o�^�܋�,!hf"S��L��H��P5%�(��~)�2�
�ۓ�	.b��Bc�| ���P`zz�^�#$���s3cՊ�@Fn�q
�)�i��Ғ[D�?<�B��o��н�}��1�BB�tq~tM��ҟ'�o|r@ܳbT�����:��:v��� 1��dN����"�C���1��cj�}���d�rzȏ�w��兴g4y��P�������B?C�)�5�Y_�|�i���UDv�;� ��/x,a(}���l��Ի=���=Y���%��?�wOKbΊ�vc�sn�ʊקiMyy�.��}�9yy�>�"M�ߌ��|�/�PT�������:�mQ�՝�!p�[��_6����ve�v����F��B���C���w��|����=�jԩ�GB1'��s3q2q�0]��L�́W��4��5]�=��*'<�{Bb���j�Uhf�V�j��x��������^��A�'��CgF�ʍ�J�ޕ'E�ߪ��K�o�7�){�W��t�����ە?�|�U���Ӌ�ʎۑw���xqg�᝗z[=�S9��-2���9����"��KQ��o��cG�>1�N����-E]��*�%�Q*�k)�IO�����������v�2����=�c~7Y;�8ur�L�Y�)xȏ��+H�����Y%����=����~�~��?ŧ]�=a�?�'޲�mkʇ�,��Hs��������K_֗B�fٝ��6gd{Wv"���\�5��*/�Xwke~Ъw�ֺa�Z<����݁��}|V��f }p�������Wǰ�~Os(���i����z��E�}6��)/aZ1�]��s���z*8�z�ڴh1;��vO0߹�N�:����\ ��o�u��Ȗ��ey��z�@0��ے�wv���v�h�bN�	$���~�R���vd]w��9���kx�����l�����9ԗ���S�n�Q!�=숐���;�Ǥ'|%N�iuZ?ȼ�5��eݝ��뾔 ����������k	!l���QՖ���9�Ի6�_X6 �'����F��K�@���0��΢���/�{�	�:��=,���?Ց������Xw�G���Op��+����)=�ϒzQ�I�y�n��ݜ��P��ofFx茧���и���r�e��|I���B"_&E�Չ�R���}f��1Uч#1	�N�
�^zn'�ji���A3X�Lϋ.V�J�)�ZF�V6��	�X��\�����l\i(u�d�����xȫ�]�8�ɮeT�$NT>l]��3xu킷�+�lϞ�3s&��nO,�mZ��R5����?��]i���1�?�}�������\�����3�>Sq�W�M��ԫ~C�C�?~�,�*w�f���ͷ�l)�[v@�`<u����g>K�|5�ܽO:�6��Z����R}A��Ā����{%�5��RP���V��'�Cc/>�O��W]E��U��zQ4��R�X�
��ia�~�l� g��I�����@�dfG��v.GZ�0��xj`�������M���/�n�.g3=�x$�Lڦ4���x�*��{��I��n)�C�tIwI�����tH�4Z:�C@@@ZA�K�C#�����}��{�q���5�̞��^k�u���Qɿ)5�Q�Mc8}`��)�F��a���8>���V6Nkj?}�d��7�|�k�+l�KX�������b���27�%����H�`:�p̷�7�I��`~_��[j���l�@�Q�����7��Ԭ8�:�_��bEXcL�p����(�՝�~������,�<�)���Y�����zJ%�E��/4J4J���/K�ϻ9?�Ç5W���8��~E|N��j���ѱ�� /*ݚ��t�%������]��A%'����,P���_v��2�T�T�pOU���,,�w��$��X�$*�R�U�>�>��;qM��9`aM��o����2�Q �����+|�b�zѤ����F�(ʎ&$��:���\��HJ����1$s�l
1E�|�_y��&Vx���I*n z�dhw-�/��� �� ��\<2��Y�5C�����xF����幰+�k������!v���璀gY��2[��)f({B�r�B�,����l9q9rD�E��]M��a]�V���εhj�.�����m�=��� �Qދ�׺���Ȕz�� ��x���PLS�p��>Kb�>+Q%�x&f��.y��<P1"�	�٪&7�Y���3{O<'���胥�}��eO��ǜo��Eշ����/��K��z�H3��2�a��ʕ,�����wV1 _dG3�YX��'��f�8R��X�'f겚��j��1C�ƒ�FW=�ˇ-�$���M-����
�f�=ha	u��ȷ���V��sMh�&Z�}WU��q�d��׏�p����1/�̃�u�m���#<Z���J��wD�`m l2sa�f��Q�/��U#�?���o�$��_�/�%��X`�M-no-�4�a� _���0���x�v�'D@P�0wx�����m6�\9߄Fq]ָ`�Xtd��Y��H�f�*Ȓ���s����c����k�Cc�-/�<D�ѓa|�鋘�iT �&��6ƀi�E�S�+7��|w������{G���R����]-K�CY�d��	^�W�`Sg���L������d'�Cf@2?�]��յϒ������kE����,7G�������r>k*���-��@�u�ĳV�@���k�������5��3�1��	�Wm*�`4J��
����fS�#E�~� ���ao)��8"�:,�X�iã�&�޵��f��^�jn�*}����3��L�f`>�%@G�ϕ���_�<�pkr�\�˳����%���B��֓�|�Ͷ�n9���Ac떃h�<B�-�~[�p1C�a� 1 o��>���Q��O�� 3d��2�E�RQk%�<|cx}$�x��WN�w�}c��A����O����Ajs��/4O��ʵ��E���IH�A��-������Q�UnȒ�� J.�2���<���6tW���k��g��~�VAN���;���7FG�x�;����+��F"i���3+��Z��0Ů�ٰ˒@By+/2��s���WE���k��VV���.�iD�BX�@q�s��yI&�w�jq-�E� :�0�� �V���oق�A)����ف��ʻ0>$��gnZ�@�h���>pZ�Ҹ�haL��/�ܒd���P��D�J9Sh�®}C�b�ƒ��k"4�k�-f=:�M?7�C���}bɜx_��Q��~������=)�bI$Ե6�R�.d�{����յ�1�W�~�%),������zpW��\�hޱi算,h��̺��y���Y>NTP�Ϫg�a ����K:� ۇi����ս7X��fLL(��Y��F,�e��{�����O�{��a��V�_���3�m�yW$�����}�����;x:���!#���d�c�W��f�lk���HPS���L�Ǩ��&Of-$����2�
���[D@�=X��;��vr�1<r1�pL^�˾޼ȃ����y3�3��:&E��6EBT�GR�'���[��-bk��L>��괅]�S\N[$�|}s��j���� ���^������fp��gH�1G%�{�J��n��kStn��,�'�U��o�g��>�� .�C�<oƨ���wh4��b����J�qR��]O��Ȝ�Q�����>A����])2�(�Q�zG�8��N����qY͆%c�j���$UIC3oc�~��O,U���p���2���˛�t%�g:�j���jҰ�߷FQ�~���/��T��
�AO�_�s��(�ns���[J��7���z ��X�J|�m�n�<Ah�V����	�켔��֘�����0�W��C�Gʟ�}W=GO<������?��M];I�OҪ	������򛰼�
`vzB{�@q�ީ4���S�G�>��H5-����4��n�K��.�$A�=���M�ɉˁ����7�l�$��8����Ai��܇�f�t�}���%��U/�U�[`/?S�U,���yH9h$\�`�\�� ��Ѵ$܂[g���)�/m1M�޽������
t�����9�}[�sa�7Q�&��^��;��!� �R��֫<|�Ӱ�уS_�TR:�b��9+�A,$���()�?Y�g�R>eM�L����
*g\u=�{9A��3q6zGv��*�Dѡ&w�m!���\�}bP�w�Ი��	`��,'r�J+�������Q�D��2��.�Z���޺�Aw��}8r�?/����;I����6+�.��΋��1uM��!��>e�d������ɸyK�Eq�
����.n��P��|sjFT������YS�8��c����m�ى���RZ�i.�IH��s^�9�?����W�9Cw�!�����$� 3"×R�%V&j�(V�C��qRdX�2��ʺ�`��%
�p�c�{�ث�N2�:�B��'�~�խ�� �I3�����c�{��}��/��ս�X19�œ�>VU&��O�M3�Ԗ�e~�?�go��-��8 �f7BA�+�sG��p���;K�jb��Z�]=�Rּ��cq2�~~�w����A6Ũ) �E��[w�Z'9;U`N5�1����f��G7�@�~x��7�$̘���#��#m���5�\��/��?�9 �zʇD����)�"ӕ'��KzZ	�C�����@��'|E�f��P7b[����+B�p�(!�d�����h���� �H�'�݊�T�FY�zh��){g5u;+$ 4T��r�OK�Y�(�n�l�ܼ�`�ѻ��y+#��17�
�c�}�
@���K��W�Ŋ��f��a҇Q��R�.r�rBd���[zƑ�&>V��F@����Gdף��v/��r5�NEGwU@���+������0mm��]U\�q�*�� � '�Y+���L�4Q��ɑ��*��p�-�o�����H��E$���o���8:���*)�٭�NV]a���(	}0J~��5���X�9)�_�h�,4+��>��K2�ͤ�+��eк��K�9U�Gd�����	�;B���c<��K-\n2��ٰP9y�ݙHԛK�-2ii�����Pφ���M��?��`��s�v%�'�~�/����I���b:`1w���w�e5_Q���pjqAд�Z9��Qēa���`��8T�����Q2C�FG�S]�-Eū���xI35:�/{�ĝ��E��q>�`N��uY�������+{���5˲e���WK�>�Â�{���/7h,�{s�A�ɂ������2��Ӯ	��J�@��쉸�<@�zL�n���H����ŭ+B�����j�ҽQ�]��B�/[�~q��7l�\�o����_ȐU���ꋖ�������Q��e
�j� ����Y��)�4!�T�J��a��뛫{[�����`/<t~Bc��rI6������N�3)�7E˕��I�S!�}�&�w�un1)�ar%	_���{bH�&�Q%�d�BNv�%���jS��L�	qr�	����.
��u+�(���^��@z��`��\r���V=�Koʿ���r��Ҡ�ԇ�ũ|��|w-�q����g.��w�m��7*�����Jh1�M�y��XR<+�¤e�t���O��!�\��?ZJ��FEf�o�̩:s�':��@����i���cUQͧ����P�_p.���X BB���Ec�B�#���bɺ}�ɓ�]ů���qO�߭c+���Ν_#�,�Ua��r @�L�Sk����j��S����.ch"���:��,������҃$���B�(�����N�!�v�oNr�b]��q)�m����(A�����%��f�%A���Q*�� F%�qs���a*��&={��`ؗ�v��p��i����OBNǝ�ng����`ҡΕ9��7��M�w�烂8ۇ_;I7-�@I?��I�4X4��A�B��$Ԃ9<�0Y���%,��R���S|R��T�-�!g�X6�����~�J���[}/�-�����At�3!М+�MN֢a�ԭ4��1��+���	�������q	#
O�d�C���ߋ�[�ye����n�ݷ"��X;Y�]��	��1YQ�i�{�C?����K-��֯[mٟ�<o��J�sp {��(vQ����a�]�+�EUFLʮ��:a8�a�hfLT��>K�A?���%�־��k���+)F�$��V J�5�z��I��t{�ؒ��^
�R����v�V�ai��U��z��Lƀ��_kU�&��2���L�YdM�̛�Ŷ��:��
�3��0=..�SaBBR.�rCei9�T�?0dְ�E2@�D�@�fdI>�g�%GIbת��0̷g��-a�$��:%0N�T�����=�U�ۼ�2�����1u���(��v�ła^���{Pu[W�'/���LL�����Բ?��Y;A6���q���$��-C7X�Ke4��0s�@H�GxODa}K��3"��{�uԟJ�,�)�V%:'ujS��L>M��Â�lj�Tݱu1��(J�U�&ۂG��B��$j���בŢ�ω3!�tӣ���14�a��߰�1�IK����c�o� W�9D��a]�00��-Hv�#-Z,���O��niӜAJ��yۋf�c{4��{ĠL��{#�ݧ��y��U�ꗫ��\��4xޯH��*`��(&���y���a8�^�"��?N���Z,�@�QΖ�I�]����Rvo��'�Yw˯���������{`��Q&�8�j�F��%EI���tYom�p�7/}���'R >?�3o�7R���f�|��}c��#bOJ��'I�q�������Vq�
���y(�0#
h��\�~y�7�C�/�e��4�~}.����P�9tQ�g���GRN��m��p��1
y��%m�X|&����Y�w�.�s0-<�7\(�݋%�$��Fߏw��wXy�l�n��>��P9%����0�e/Y�.z�����Lm�&��>�#-�W�40�g�!�rǯ��)4o�����kxW�~h�_���)�"��L�)�b��E��t��B���ޱ������2k||�L%`�ඹٽ��e���c�<V�	u���O�[��.{�5:.G��X�s�C�Q=W'~�B�z���e�N�xS\�~�	��_�n�}$oa��:z��{��E��/4�|۽\~�4�S	�35`��bl%��{K2gƳ���F~����r���;	��?#>�����p@d�`�$ò�TX�R��t�b���.fA��d���vic���K�F�s���
'�d���u."�'O��ML�+do�e+tFi !�JYr�U�{
���
��	��)����T�a���ڇ﫮Z	3K��赓�x�G#��8ykŇsP�|�w�tR��g�Yގ=H����\�q���ګh�
��#1��j��\�n
k���S���g*�4'�]p.�h���6��,y�g�d��($'��6}��^8�Y\X�|��V�Q?�@����3�Y$`�[���p[v8ܴsC�j? #]�yg��d��*sv���B&�p��X;p <?W���¿�}�$���i�]`>Ů��j00������r�9���{��:��/��}"�S�,��u&�z��n�2KV�"@��2KlL$���#_ۡ�^+)4ݾ�cY�Op�~��KKp.�Sǝ��C��`�����{����ġ�y`nUnǹ�5*��#),%�T�9/�";�?���0O���u|�.�*��|���:���~3iVG6��o�l3��)����}x��4!�@�Y}���]3��9�٣�ѩ��I���ԑ�W��b���0K�gw�ʍ��F��P�]O#�����[�~�~XC2����u�x�	����Ñ�w/�=5�����;����j�U�~N��4��a:h�(�|�Ǌd�܆�������e�5	�`��3�׎V��x�E>RI�;�G��9���ԙ��'�ۊo�dN�|bm��A?VF�Yl��[-�v"z��ˬ����<f\ F�%��N�)�Ů��3'��ިKuL�S�#���)k��0ZRPw��i�UovX���N��uB>����0�3:�7:�	����n��f~�m�F����j�M���`ӓ
q�INH�"�������1���N$?-�XYM��3U-R�;5+�#�.}�&��cL]����f�����:�C�o`5����qTj��L̖ڽ���N�^=DV��.Ol?\�Ҕ�ݷ�1��������� �G�����$v����ߎ0��3�p��{�pK��XM����B��"6�����֑��ۃ6zh}+ib�������J}�'_�*�+�no�<�蠁XHˑ�P�G�'F�1l�ZKH��$��Rn�i��x�#8x%���C�F
x����L��=Ut�7�YqQ��e�oL��p��h�j���f��ˆf���]{�$@=��P�I�'DI�ǣU�q$0,����D܈��s�Y��ɴLi�+�ܯ���:����Ϧd�Ur�~'Nhu��)�����`�jOQ�
'X���1�l�t+j� �U���!Ro�_=�(��h;P^���AvTܑ��G3>+�8tcj���e �B~nL�V.���9�AŞ�rF��WP\�ٶG���T�r�Xb˪��{�"��	x֤Q{P��2�C��&��p	-O�Տ��vk����Dr�wq�c�s�)};�: c%+_>��D��+�0m?Z���s��x��¡�������8�34ՕKw����N�!���r'�tܮ�ZXqWZ��M�n�Ϭ��[Ph�[��D������ПV�K��[Y7�~qZx����س{^���W���:��&ϗ��|��n�)X&�z�)1<pt�G�^�U��;�i�+�t}���0gF0�%Og�)I�6/��N�'�q���MLftg��eU�W�,p8�Ш�~:x�2[�����v�Vn%��7�dP��FRE�}}򲡐:���n�¯#�"��\d�Q����-�e -�u&�_�( e��4�|j�O�lU@��~�Xo�:���ک=j���mm��&��
f[_��֍JP?�8eifp�9�cA�fp��B�&���~Ɔ��)�&�z^�TZ{���X�Y�ņ�#O�#gn����L\��K����ӻ��V����dyܽws�&G���p��V���)�\^�<*�)��B�E�J�k�H����Jٯdo�y�L�33�Q�ṿՅ���d�Uapj:7� ��0̼�j�r�Z�[W1��!㌒1��2��\c��V�R��mp���u��n;�T�]!��
>ܣ��N��� ��|�r�^LU�ϙ�U�
�;���u��1oo�#V��4��y[�}��G���������?![�2z/�.�$䑣���&���8�Z�����su;�x:�s���h��nK����d��x�({>:�n��\����A�z��P';�Ƙy����M�_�"co��VEE��gF@��%104� �6mSy�\xGj�c��ۆn�¹7�������+�!V�Jѳ΍��_>`[�ұ��F%]�i� �ٴ��͑�3C�$��B�/`�<�Mx�� �ۻ��ߌ�f�r����^�R�S��4������b��j�b��=��.��t��5B������i__H�q8}ivdtj�{�J�$3�J����P�7���>9愃��s�q����z���>+�ywcX�W��dV�����I/�w�E�Q�_6����qF���"S�,P�_ۀ֗�7i��b?�b8U�1e�L��uq2�1�]h%a�уa�Fn��,��n�3��6:��#�frƢ������1d�X=rȮ$��_,xm
��\�<��֟�$k&4��G�l $�f��c�H���c0�IN��K�0".;@���d4�wW�{���㊟h�判��F:����6��ar�ϭ�sS�/3������0~�����xs�+'�U�}��-k������Q�a�����"��⠙l[�V"���J�f3c�l��س+����>�-�����f�>��B�^ 7�!zqyȑ���%��\������-fi+���:׼?7�Xh�s�0�;a�u����/��s9����LP��o%MN|ҙ�}�z�&���lTp�9X�Y}���g�T�b��DWͶsN�i���6|���|uޱ�i�Z����Q�����X�����.Cެ1Hl�b�lB����s�y�l������g�����7�t��&�
��\�$U$ u�p�b�;��n��>%�t]�TC�. I����zJ�1u���K�8�ޠ-�AA��xpX���m(ѡ�`q2-e���I{�,0��&��a�ۡ�(5���!d0G��E��(A�V�0��+�&�!2	vC-J}��.@�=����f<�<��`���A��BËw^p�[ae-�gAޡR}��8�S���]^��t˦݂#�$�FMc��B�/��|�}�H��a
�ǤK��hdou��N׹N�6T/��ED���'����_E�f�����aU6�V
�z��%�Q9�-����8���Pb��
1��&mX�����.�����SX�X��r�B���q���)ä�|������d3��V�Jt�L������pW���] �8�%&���A4C�SEu�f��QF:Xť��]��4$k�]潅!�8Hn��{�}��)��Y�r�p�A� ����8��FJ����P�~��#[ۯ);@�c.0Ƭ�`U^2U�g3ûu���4�֍ft�Kc'�Fj�X�<�qq�?��}~���&�Ԇ|BO�fU���&s�g\˷H/�v9�F���1}�U�ɳI��s۷#�z�qT6v�6��lQ�kr�"C >�}�\�'�9��������w�F߇h���"]�� ݓ`�T��WHMoNUj���gi���ͷӄ3����_����l)��)�a�ԡy�/(Tn\	Uf� Y���!�ľ`����K���Ej�+R�Ϝ�����:XoU���P���*ڲ�x(�e؋��� �u�s���%� ��<6��d����B�W�ު]q��f��&c[�9��n�{E���%���.�͓��v�����@�[��:,�oJQ.���k'��Q3:�Z +�'�F?[�#l�˱��|�d!�`d��)��ؑ�I��m�Ǖ�3b�B����H$x3-Hv�F�?@^A�nG�=7�e����#�*[����'2�����W1V��$�7�%��r�G,0Q��8���E��*����`i&Z�0Ӻ�ʌg�~�2�$�a(���Cl7�� w��H4nX� 9,�<␛fS����yQ������?sJw��f�'(���qo��O���tG��U�&y"n�g�:�B��(܄7Z���l����NPM^.�2�����_��/A5�����#�.DK=l�"'4�T��a��n�I!X�3{VCe�/=xKN���J�KIl1���r���[�	%��'�푫��͐T���N��?���xS�� J�絊�f�-�X�]�����9�e+���Z��A�V�Y��A�q4D|�So�Y�w����-rV���������v��u���D�2��ܙ:��A���7#e�'_|!pο��`)ˈd����6P^&��ss����Rk*[�,2F-�QO�'��	�L�Q�3 )t3&�w{=v�S��}�02b�'���+=;vO�v�}�w=�!�rIR���  �Bj՛+��m��L���}���\�4�1z����<����q�}_�$�~��2%��]��I(Oi��F��������ʹ3���t����$�%&QA`�K��ǿ��%�p0�η�w`�9�ӥʍ^
���lE*�q����,�Om�X�U��y�J�J��_���$�.Ps���r#r��2eG��8ϼ2TR�w�3k'��|��`�L�3�R��ׯ��r�Q��W^6���	yߗ�)Ⱥ�5۲�t�$���`��@Ԡ\JmsU���L��h�\�Ԙ���������u���;q��6�P/���HfY.��?�1�2d��s�"��@d0Zr箽W��L���%�~�����@o�{�o_�N$�~�U]_>aKu�?*���^�0 �l�u@��@�Ƙ!�ϻ�=�w@�
J�Yv�4R���9�.��`����W�F�W6�������ލ�x�*>>đ:�Cb���E�pw������˿	�
:���Z��!TOc;�k˟g���1{2_o"{��	�j|�pM�Q�z�+#Mߡ�Ō	�n�0�yGF�q�u ���t�Q���T�*#��$Kn��9A�;��O�zc��с����zJ�}C����2yed���/�0�G�ꡌ3��$����b���n��ꠜ<����V�C��B�i-{�i��vV�di��fz�/-4��3��hK��j'%��m�;���'1��q�", �w�Ma��={D\]P!1����?ӭ7���h��Ԓ<d1QNR����
H<��Ё$ᵸ"�F���p�O���ɇ��	� 7��\�sE����>n��,Cn���"B�hx����+%���� @����8Z�\S�Z٨}�a�\~��-���,�_���M8�heCӯ
������l�:�e��[�u���x���^tSv1�"��� t�K>��+��Β`�y�M�=��Zo�ț36����Dþ�O��l���@�����=N��
@��(�t��i�|�ni+8i΀�cl�H�-�}���3+�:� )<�g�_=�[��wiȷ3� 5�T���9a4��S�FW� ���tH���bt��S�&bP�)�i�9�;H@�~�S�\���d�f33��`
��l�[;��=�M������Z���[M:��S�!���,�^�{#b�tڦ�m��Eƞ��{��JP����<��<j5^��Uf�g7 $P���q��%  �$�ڥ�ʤ��Saw����w91n�uX���Ư��V��M��*�'͓�b�o�RW�h�J]���no���q���^��q�0q�H��'Ǳ��z�N�g9ӧ!jW�a?�A��3�d�s&�;J����Fh�����U��O��w�yuuS�md�=�ޑ(�i^;Q�#�Ḡ"O#��b	])�]�%��(ZpT��d�R�d�l�/M�#yOni��
2�ѦOߔ���	�!1k���=��;�+�v� ��ĥ��{�q�A������{,D��[&�d�5��3Q#VӐ1���2Ht�&�H��*��@e����h���A����`�($�Y|�Ǯ}��Qd¨߄�h�RqۿӽOu�T�N���~ w��_�,>��z�~��B�v.BݮO�k��y��T��C)zBk���X
v�q�C������e������LFM�ξ�\|�oR�Wi�����<(�U�K�5[t���Nͩ�sQE&�X�������թ�
�
;i����i��|�c����(�O�܂�sF/�*_���Z}��ϱɄ	���5��&I��O����(ѹ u����w���??\�Eذ��y�ٴ����;���`ȼ|�r: G{Aip�a�7��7r8W����(FP��]g-g)c3UE���Ìe�?�o0��ij_ �M`�ԏU�o7��KJ 9
��I	V�Q{w���Al�#f*Aqc�m/Yi�,cߗʠ����<Y�х��%�τه�!�_�����UK�"UJq[���nOLC/����Q+����sF�T���"�R��e�k��ȧ�)��FNzblܘA=��z�Ne�%�ZY��6>T��v�sp�Qwi���&��q$;I�@w-�\Q�D����s��4�o�����(|�|`���³�h ֗�*V��l���:��-���Uٲ��|ڗח4@��?|��1i�6{�;�v�e�
MG5����%�| o�Z[��\ڗU;�vh��B@A��T;n�yy��-`��$��B��.O�&C.�Z���=�^ N<9km��m��M�ܲ���I�%��)܍�f"1$�1@i=>Fy�[gq��uǾ���<6�n�|�� W���r�/�l��'ǀV�M��h�D�X� {`�à���<q�x�k^�%�j�W�0�I����x-1������O��ׁbM�� Y�{���1�PM �c0e��<db჈�*.K��U�%��.�a��ў`Y��)�]�_zх�w	G�6L���ك��3��2�svD�%H��g�1؎���~��؍���y󤇸��p��V�ϻ{TC+�r����"
C�H��^��y~������FW�L�����9����0F���9(DJs������&*J&��7A,��w$H�]��7�k�;�u���>�=���S�#�d	���P2��,�-�l̨�w���lM�Vn��Y}��^lՐI���}f�V�v�U{|�-���R���3L�,�����ZEvr�x�[���I+�Fl+P��j��_�(gK81��1,��<Tn�_Z���x1���W�����ʚA���)+}�&�z��M���A_]�<$�2�����Gq����x��ӱ��~�G�
Y<�Z�5����).��R�Rf�^��̓��qn����ت����&�t`�%�s�w�o����Q=���(��a�u�;�,�8�VX7~낭� ��u!ՀX�K�����N�z �Ե��?�QE.(U��B�|O�~���[@i�Ѿo� �D�Ϛ�0�7W~�87�=��m�j�l���!x���������[�������~q;��V �S�bn�O�m�M�;�w�O00q�0�.��v��oTۡ�X���|�ڜ���J�w�z�
+�+��'�[���������J��}>�T�n��^�$�^�~��f�`��m�Ɛ�d$5�j��K��9%�E&�Wl��l`r-+�dSr�^
�7�����|!�mZo�>er�o
������t��@�J��re�<�J(Ҥ�a����<y�E��4���*PV�z�݅�-�I� &��7^5_�a�-®�[�9��������C�7rv�����ۚj��N��l�GC_�����ؐ.����w��ho��
"@< ���_�2&�n��{�d4&/�����(a(6�Zn��j��i���Q� {r�D��1��
��Ǫ`a�+Ć^.����nR�?L��v.q{U�a"�ф@tL]����Z�:;box�����BN:����w7l�-��H���e���l�c@�*y�|�T�Ǜ	��r�ҷ���I!��|����2ʘ�d��q+���&����df�m�x4�3�u,��c�V���wms��f&�lk !oo�t��Agg��O���`��v�-7���vk��2����9��K�l�V��������͔�`#D��1��b�Q.�T�7Z睱x߈�����co��	F�/�m/&yG���|}��&S�UF��f�����Ɓ��/�I1��s���!�l�Vi,Ș|(������X�+x*zS¢O�"��*Μ��`���$���dg2^�N�^��Ρ#+�� �1����~x5^�*�<(��&TNsXy *�P���/	�\.�T������,Z@�n{S�.'(�Y8ٞ�>ˌ�Wa̧�]���=.�6�7�k�!'PF�L +Jc��i���ٴ[�����(I��5W��3f�]����o�)�T�w��so�".J"����Z����#4C�V����VV�V7��� x> �"�Gn#Zl0�9;�[d��sO�78�:s���g"nP�Ŕ�E������x9�-s@��&#ŝ�p-�;>Y\r��1l{�-[�BU&���w�=A���kW�/ʀ�9��I{���騢41���wi�;��,!N%�����k�?���qZ_�6@���b݋h�y�霺�W�ga Q _}[5��f�����<���k#X%��eivh&6��ڡF�㡝�����g^����925 X�χ�3��s\��"�6�y����l��,Y�Wl����8��㛞�-KB���[�V�u��ko�*�P	��Cdo�8G�gL=�����$�ڽ��Ư"W����G�`,�g�k�JG�츕�����CY�(�e���}��D*q��$��#;�{�vT����^K�L�Zo5�XJP������L��1������G��]'S�wק�x� a��F�F�1fH���a�A-����{T�m�WyY���ޓ���W?h��mö��G���c4P�Wo��&j�󋤇�>�Hs�Fe|�ٛD"�'chn�RX_�3�v��q'}�-E�Õ����O�Dd?�G�d���g���P�驨��
���@/��B,�:�f���1���$2�����t�]À����d������0����A�7�'����*�6���m�{!����Ǭ$z!%1o�rN3Oޗ=tU0Y��K��`#����L�_Qwp����F���d` y���@����'�
lQ�����?j�?�=�x��Ć]�SKbqV��nt����Z���aV�J��Mbi5��$��r�tc�v�X*>���M���қ�Ӕ��aS�V� z���P�XB��8!Ϊ�لČ�*S�i���������i�F�����RTpLU��k��T���1�B��8?��|�GG��r�2���'3�F��b���w��ëD�$�;(
����"�a7'�j�S�W�pӓ�6�a�!�6�b潦w�&��}#��/�32�#A����b-��&6��p1�����:��������{��,�Y���1v��a��/�����������~�͟ѳ�{1��}�朢�b��K����%]�J�aG�C٧��aa��E��;OAR�#ޘ�ρ��X����s �H	\�ܠ�/����y�tg!�:E��}crfo���|�]�m��#��O���Bҽ4p��z{q��M�&�+7�g�����p��%��<��& ͜�P%v�ʯbC�W�辛	$ Ԟ��5V��[��f��,�;�)셛�G	�Ƃ.�[���7T��2ެsM<�y�����o�ܡ�$���PX�hk�M��_z�޲��}�Q���ݏ�b�aw��*�ȭ|\��u�x�2��X�kAj>z(|9��ݼ`�;���.V���������2�\�R7�
���L��GYl��}dW��1�*H A���5k}/ ���G�]z��g�ܜ��F��y�����ŗ�M8n�����[9����W�a��B�ŧYZ�il��k�k;�e6�2�ǔ��j�tYϦ�z��l����i3���|�9��v���[��zYc��K-���PHk4Cʳ����t���a�4�%weRjSZ"K�e�ǟK$��Q�Ei�����|?:Ǵ&<JRa��;z�9��h��euR�St��:�Ն�cM֠�?|�s�ܧc��9+�Չ��b��EV���G�Q�d&�w����d5,M�U�{;<���=��$Pg���3��
����4��� �!��٭[���kl5�U��H���!�)}Q�'Ś�#���ܜ������	1�[�+����O�����a�"��+��럯|<����/)�Ԅt�H��~��m{��B4�7�bq�� �cX���(�b�6��*XI������YuY�q��� ���3[M
�w�ʍG�wi%ܥtdx!�^{V'�N]��L���C&�ȋ���O�j�raЧ�$��無�IU�,A(dz���;6�J[���j
��c%-���E��lgG����(	����e��u��EڈSR1���Z?��c�¡9k�p�mȣ�V�.ʐ����)��ϗ�/����I�4��A�i*p�J?*����
�x%��]��}��9_��!�.�<�^)��ݦ�E�_���8����~��|
�hg=����y
⇉6�H�"Y�+��P���]e�Im0�[V�0>�}>���)���J���w
�쨪�X=����B��,���XI�p�A����������у�����Bɓ���L�aBr�bV�}"�>7!�֑'Q<"�k������zɪ���o�F#�[���>M}H)��=�T�F[j�
����T3�d2S)0Z5U����~̂����Z�o�9�!��f3NxZ�}���k�:�+ [�������Z�O�P�Xy��gz�?��}CEe�y��0y��K��ƑT��K�r���kIpLC���CZ��.�A�����/����񌼵�к��5-)fq��S�Rq4Lm6̓�Ῠ�8�����U��T�O~����/�oBQ@Z�a6SN�<�E��\����X���wR��
���O��}�W����ĸ�:J\`h�d � ��\c�=��(/Q4�졈w�I�H�US�������M[��*�@���ߣ��Ot�]���Z��M2R'����M��aY�H3+�G�
Yn�9F�4�����5Q 3����?����݉U.+"KǇa3�F�%�-F��MQR"\[EȂ8(6/5��w��%*���ը��ÿ�M3����g��d�����^�'k�ȁ�q���F�79��t|����9���"��<�{�&��K�<!Q2DP��G+�Yk�ۏ���̝�������ܘ�@��Om
�p:�j��ދpP�g��d]r����$T�e��s�i�ɼ���k�Tp�D�̟�����M���'��a�7*����@�X�-��=xa�G����璎����2��/������=�6UǴ@G��!�.?�0��C���y�8��MS:�d��cf�n���������M�C{�����>K�[�V#aS�|ҩ+>J7��i�=�3�I��a�;Z�CL�ۃ}����[�k���~��x�<}u@T��5!!� �4*�һ��H���(   ���!  �tIKJH#-��K�RRK-�������ޙ;O�眹s���At\ta����2]����;�΀e�T�G�;YJ��J�JJ���Y*�+������IU�~�����Ef�� o$H_At�T�Qi��߳���703@�<�+�����f�]��G��ז+-:���$��Geɍ��^��^�M>�����e��SOq�]i͡���-R�@R�t쑘>��R�Ⱦ�g�ﰒ�B�.�����Ѕ�ӂ'��( A��Rb�B�G[���plgѺ)�q�/#�M����5���:��h�Ѧ@��BD6esa��]`I���"-c6�������H��G�N�s{'>�:���`VD�r=t���|	\�O��������ʭ�#���Q�گ27�zv�����;����v��sky��dY�u�l��D�����w�G�gj���*4cv][a,*S�w0�G�o6X]#d�����>��إ=2,+3�u4���kp�����:�V�m�oxG�;kKf�� ww�EX��@�p�;09���Gq�>Ů���{�҄���r
�t�oa��� ��+����`*��g��@�0�O��!��o�%f8�D��w���;8���M9j9���Y蚂�V��]��<��X?��)��H���sY�ٞ��nUԧ���k�1ή �B����<���@�����\�Q���<"��5�X_9�H@t�>������bo|���dZ��{�Ϙ(l�J���?ٕ*X���?��������q����y<8�WDG)���lmav�ኂ�]��`�88ֈ��ޜ�ƈq���f6'NkB�p�m�F,���?u�#�ĕe���N���6�kE9&��9�p(�f' ��]�=M/��Ƒ-$�K5iG����K�՞
���&pX�C��Z��y���d	/�gE�͸K�g��_%NNʕ��T)%�هu!�i�Yf��ʪ�"���X����o}�IVGN��Y���趩'�yQn3cg��`���d;X��#(� �jXxj�(V��	�74O[LWO��.;�Ä{~�q��c�G�G�KՆ���GnGn��?�ƌp5����&�Higo~Ix�Y��f
��[
`k�c��KUwY���}�*u�#a8q;.7~��5MG�|57�ф7c�+�%�Ӛ�����/�:Nv̘���d��gcp�X�x�>t�P�˓gǒ���瀤M�u@�pX�+�596�!��&�4w�7�X㭜�����]��
�(�l��H�+��>�̯����H
���xI����!�L3Og!M�`�^I�����|��J��`��koᇰI/��v.l�B��$�K^]=�<\Ύ,Usud���T(��UF�^���$yL�*��i?�����݁/���o���]~�B�8�M|0B�A2���SN'�����.����U�-�+~���GkB�%6q�0]�5�SΌD���Ӌ��=�Y��?�&�)�2��	�O`�1:�[���$�*=\�8��7�ې��H���(^���ƹ��8#|���'"�+o4-�{���zUN.���,����^��B�6K��+~|ы�ಂ��
��
eK�?Hc)�Cr���]�z=�9.c���i��V�����C�x�*QlULmܐ�ҫi���]�V�m�M��*�����dcnc�;�A�B.__C7�� �4��V�1��:�-�� ���;��w>�7�Qڼx�^��O*x�C̱}G�u)�]�^���ϑbWZF�)`����3#L�Q.���3��F�˿"�{�e�3����%W�
�ͅ���27�3�����/Ё�~T٦�o	�d���A�H���y^��j��K5�::�chZ�oN��E5%eb���%� �xݜ&��[z�y�u���N�:�:��97��x�1�頉�R4��8g�AIcD��wT�0_�a\�<�������Q蚝����{��E�����Q�{���7��}����,)���_Fo��^���~p��^�R��5�����Fq��Q�ݯ����ϊ`��m�͂K�mo�csTK�M����uw���ݲ���?�00(�aO���:w>n�: ���R�ƋRu�94⩂\r�����Zɒu�F۪��
������{���bk�$;#2�wm�&G����P���ōoۿ@�u�ɉ��;tv��/{v�������:B��]���[�U�z.���i{���"�������,JS����FZ�wm����z����^�]�D�?ֹ��cdj�Ϳ���;1������+��| �V���,FQM��o�����$��;�:��P��n��ݷ�R���L��
v�h[5�O�:���O��gw�S����'+�:%�w:�$#_{>~9��6�P�<�s�\ii�G㔴��Eɛ��hD7?�:ι����*�����1�]M� t���b���ie�-Yuv�t>�Q<?\�	fƵ��Y�<�v��e�����'D���+~����;Gb����r�N��{���z�pT�Ik�?Sk�^�PC�\-OM�3lP��xQQ)i��c�e����7W��Vfe����<�KZ��N���`Y���tI6`���hs`8t�p��nE|}�����G�ǷՀ��*;k�h�o3_�R"ھB�fe��=�f�"O�s<:�|J*�ԘQ���9on�ߖ�"�U��[�rX�>A��kk�~)��$:D��3FT�����&kg>;=��fl��j�RX���-��ک�@��?��8CUGD0an�XM���/mα�kj���4K����{��������_�0��<`��ժ��9*:U�v���/T��������}���@u�_H�A���{r��?�@�7f/ϵ��^��Xޕf$B]�Cɹ�������xB�a��P�@lZ���~u�B�i�ew�P�6�u��R�
͵9^c#�(��dr-f������,��#FBc�x@�*��%|i��O���]�{�A�fS'G~()/��^� ��X9R���-%��$�Z<��|� ����`ΚD �Hj=θ��4򨴌bGYqo�$[H��at�:��v&��E�ٶ��|�����ݰ	�q�z=9�ƒ�!��II���]�=W�#����^\>��@;��k��zzVVxZ�
s�41����p����6�������b�]���S��F5�^xKX'\�ǟ�/�uĈ�������F�ܥl�"���+U�1G��)a�U~��܇�V��7=����M���5$��'2����`���ޢSC]�+�#�nE�H���-������]�@����J�p������5k%Κ�맼�(��_!>�ۓAKo�ņVI4�O��N�g��U3�y���;�W�%�:�}6L��VS��7,��|��6L'�;Q�}���fW �!�Ф�s�M���%dIle��F���IZSy{C�]�R�I�T&��x?{i�j�냛5���V%�<���|��n�}��	~���*�c0ɲ𘇁�6y)m��l*C���~7��s����DCF]�':���0}a�2�����[�����3�2��1t:K�3�s���.ŰIHm;��׺�ru���jk���[�8p�f܂���Ǆq7K��
��)��Al�1�=���\˾��P32F>0��]�	c#&����({�V*i��qӇg��hdm@?�˟����0!�=x��7�B�p���wicM��j��qMpý�ǹWj�MS6H��+P����V���������1�7�����\�սB�ZH�2��vU��#�O������m�4>��1��8rnY�����,���c.%�c��a%�[��Q��Wu>���V~�1o��@��`��w��.<����m��_a�2��k1"O��Y�LIA'�54)f�ȼ�ߥu�L���ه*r��!�8��8K�7��}2����(m�(!A7x'�	ej ��~	_:����ݦ+U�eh]�B��Y�r����S�7��>�	��Q���	ſ�[��enV��Ԗ���?�ܻ>T�ך�]��i�}5��֟���dSL�o�c#?�bF*-M�.R����(�:o�Ӿs�Z?8�l�L�+B��4�l���J]�~2Ag�)������Nt��d�%(�EZ�.�������F�_q��(�v O=���#���(:YJ����^������V!h�����0�}7�e�3����!�y����D��Ɏ��	��0���S�����;����$��"�������i��')��=rh�楜�@[T�L��Lf�{g�[i�r-%p_�Q�-��ӯRu%iG}PϺ@���T���'�7{��n����T��|���>��`��nIU��ϗ�H�)U\N���U�����X�?h^ ��뻭�T4D�5 Tʽ��)�ܓ!X��-��A߽~�_��� ��y#�fd���W-��[&E����o�a�ƥ�S@�=0;Ǭ���Y(!�C\
&��b~��9:�s���+��#8�"��6��o�:z+Ǎ��y���MÌ#@]oz<
� '�YK�D���'�q�d�ځY�-Y�J!.A��૊*~�uYZ����d���\�nk=����E�\|oj�����}5���?bӧ�ĕ��ޡ_Sbl�]�����LtY��h�S���x-<e�(Cĝ��ʴ�V������f?��=Wq.ZH�@�(�ǥ�
��O\I��A�;��o��%�������h�ϝ�h�u;tz3��<U�h<�CQ),En]X)%��{2�.��C�Y,=���㚀�����:�n�?u�3�����+9�]�s�U�_b���/�p{��s�b�9N��5@2��_���ӓ���BT������:� �׹����B�n�H�K�R5�|�[N��;���g[�E�{�v'��\�߈����L�j��ǖ}S��t19�^�~�/G�O������+ھ���#�=U=*���5% g7y6���/뫿�>i ����Eg��IZ���A^y%��vͫg��1�e �$gl����S�r��~e��仉w��o�e�R���@��!!hlF�-<I'Jk|��k���Y+��1lq+�u��<�?|yn���vE�=M���u8�/��˳W��i�dVtД��:Ͽ����w�d�8Y��)��y@_`[�x�gn���h̫�Z{Ŷ��j��+r���O�|q�	5~G�;�_*�����}�wE�T���\���������!�5#A��Ak�n��w^�O�x���	4|��`m��Q5膷�X��888�3Y()�G����59�I	��ڍ�E�I�TwP���n^5��}�fm��ٟ�� �Nٌ1	��3��T�yA��Q��-04p߷e����qo�:;µ/,/C��R7�=�+�T~�?�Y�.Ua���Ly���k8O�9���LVB��2��w�jL:({�A��R��"0�#\A�a�E��[�a�8?�^�e|�B�N��,��ԭ=
��!I���ŗVt�}������~��ޱ�K;�&G�!S8Y'O����]�~?IDa�sp�H�mP���Xg˞
vߓM����|��B++�y�a��c�,����W��Ã�M�	���jZ�����2���.���ͽ#���79���>�{�x��~����I�l؋R�?fOA�d.��
�$K���/0���!y%�F�l�.<��3�ƾ˯$h��Nv�G�f=�'|;�] Z �ĸ0�۽Y����L^�\���=�񱾰��l=�񀜅��vĬ���}wH�x���%2��q�8��6tjVB��G��
D�� '֙	0�}V�P�~ԡ�=�Epd[��~�.���;n���V��o,_��f�I}�w:SC|�qy[�ړR)	@W)�u����O��͸�B
H�6 �ѽ>k	��O��̑Q������&��q�J  <F�+X�y��E8MWi0�����t�ܖ>�#7�̐��L�������+A}q �+�s��5,E���,��k���ap�x��J��}͍֒�����������4��ܒ�6$v@	��t�y�}N+�N���u�u-�[N�=D�FŘK��Bs�����]?`���Z�q?l)Q������@6'C�H����
�\B�j�?����ݎ�Z��d�/W�U]��И�~�9�13:H�_����Ώ�#�T�g`���,������M�x_��?�Y!�7}Ccq���"��u�����!�i���ԃ\˷�p��M�l�T��V`�5�˸}}�~��V��?��ICȊH'Xf�n@d�|���1���BK��Z A^�]էcj�&����Z��Z�����t�z�� �e��T�7�<;��.=��̚�έpB�̉��o��j�Gܺ��V'���__�n�&?��Qdu�لِ+���-Q�����eC���>�}�+����Ä9�#y�B�Ŝ�u�+�"X��J_jx�S��}�q́�W=�����nv��L�ɼ|U��-e����)�Q���Z�ñl�!F �lH���Wyv,��21L?����(q2�<���W�2�2�QK��lZ ��=�Z��(����; ���PD���.s!�4x��jw�ޜ�!Eq1��*r���ʪ�k������c�&�0Jl,�(��o#y	I:^���g��Tu�O���N��z¦^ȰT������499[k�)e�x.h��ƿ��@+��4,�J����P.�>�F� � �{֮���s^U����O?iV�H������Pꛛ����ͮ[�];Njw����&��	A��$�}0J�	p+=e:�1�/c���1-�E?��85���\@�G�:g�Op�;�rp��Kx�6/L�������V�~wR-�9�{��I���n�'!vA;H� �1�L��Hi߼�1��.�ƾI�!�o�~���*{���1teboj>W������J�dYM���JBE�I�R8�Ul���;�����^�zl���f%��'��7�S���i�z���ZͰ��]#LBh��u{���br�,=�V�.ޔd�[�}�ie��sz�A?���!�Y^e�cq��O9��t1X����`h��iȳ���/s5��2ԠD
�;�\s�������$O����v%�5#��P�?/� �#���d�IR��?³~�ՠ׺�[<�|x�N$�ɛi�OB��
�U
*-���E��H��Fqj�i��ޭ�Q�˹unF3�h��߳�r�g�$�� ��uy>�&f�L,;Z��ML^���5��&8�z��]���@�W��_�r�׸4ΨiJ馠	��j`��e�����"���k�-���[�={�j�3Ph��C�
��K���˴��t��WT�=d�`yդ��P��!��S�I��>Dz%&t�;��f��|��Ǒ2���y �9RHc`[���E���q�d�\��?�p�C_�����o��� �-\�k����s=7�q4�&U9Sd�mUB!�t�ԭP�_�p��l�m���!��S0t�%��,��kE�s��ɡ����xl*P��G�O<�1V����j)*�v��|;�͗�W���Rcv���T4i�r���U�o��9��3���w$\��chSVWFUm�-��Ǌ��WqD7|ߚveF���h�҃="�����-���!ka���*Ѥ3%��&���{�G
�{�<������FH��(%0��L'��d笽���ж�8��i�m���ߊ��)�%�i������s���h�vk���91�X1X��A��{sd�
˧��R`k���<U-��r��^Q1Wv]^(s���3��g�^���Y�[7��I�|���K�,b^{��Av�/�O7��%ΝM1L�s�7��&趓�iBAG�ť��77"#h|�����"V��g�=�c��+�n6v�^q)��ϥ�.Du}���E�乳�����������$������6��M�6~��Be��aQ�xϷ�=����D���_��g��������1*�Ș�"DG�(0T-D�
��z�Ԯ|++o�x�c{dS����,��4a�T��s-��]cCJ������mz��R]RG=�.Y����)�c�߫ç]O�~fX"�|�}ZZ�'�%m���
�d�,B����ш�؜��86S}=����z�.��c&��P�����z���2'F$"U�_��[Fu����������:�s��0�۴z	_�W3�]ёv�+9�|�ܞA��~�Ҙ�{��9s�*�'ߧ�_�����5��.o?� �Bl�m��g4�}�32G
��/�?؇;��+�O�$�L%%$���=3�ʔｴ����&]�۰2��:�cMk�7ӣ��e�����R�eʅ��I���]n���Z
S�%��#�'�;��E�+�������;�ukP��X��&�7�SB�)�����$�2W�.��H�܋f!����q�O���Y��z毼� &Df���f�60�A�j��\F����Zv��^��wƮZQO��/e��SkZx������G#���/���B��k�g���ֹ�Cۥ���ʺ��>�f������X^���5!g������Bfa�mu�Y]z�h�Qi�	Z%�_���E �4'1� �
r:��ߨ�s䘥n�VB���hz����p!]��d�>��ݖVE������v-����T�~QiU�������m��h���������:�ey��98����f!����m��R�^8�1��7 �4&��r����.�0r��y�Dl�3?��P5����fzNF�-�`B'�˧���G�(��;`�<�-��2�`���ܠ*qA���}90U�qⒶ��Do̾���B�g��
�%v��dN
:ܓ{�V��ӛ��ǚv?���6C���e#8���\��/A���}�9	>�dh�G�ڝF�܏�$?�/����Dh2�ק�����`f�����D�8��Ҙ�p�Y� x�Ϣ��Q�+����,;炵�\߸�z\+����d��2*H�\|w�\"OJ{}� ��3~��[���BM�����h�ŸRl��3	(���	F�;����y���Znl�Pz�	��ʐ?�	��Q�I$�@��?�����ج�~Qw��	�ݚT��ia������(X���1�-ׇ��O���pw���ak*��9��Dy��,!f��������nA�,��5�O�ۡ]4ۥ��J`-=�G��i�RBа��貹�ԍP�f�$��U��"r��=�bﰡ!o����ſ.A�,�~_萛A� X5��!:͟�(4/��#MH���ʧ�S(�1C|PW��˗�$5��p�+��iSn
h�R L'"E�	�TZ*h��1�d��z���»�Iŉ�˩d�4-	���4�$ϲ� ��/�
�Å��LR�-��|^>�}�㯂�^q�N'�L�i���r ����9Bv_o��X4��$�.�Ca��V�g�f]���b�L��!L}���*��\N�rw�v'�h��r��A����._w��:���@���Q;�	>Ɗ ���� ǅ.����P�36^�"D��y��i�F� }�����n^y�8m}�Aʖ��
�C³�SO����wSi ��}��J������|���Ka�hQ�>Dſ�\"c�`�/�Q�j�7�H�[a�ܕ�z�췗�q���B^zH��1}�13J����:?��_<�Ji�K�y
�j� ��7�s�*vg�>��G!��sQR��!tP�Rӷj٩�׾�Z?������ +Bpa�Z��[*C��9�<���( ��)3-\ "�W��-����S���쪏OD��@��L�Q�����]��Xr'�ފ�H�C����Иi]:]�B����k��!w��$�V*�Kw�7.�-�.����m�����8��=�:n3�����B9 ��?��=�H��ؕ`mKh:����.�e|�J�W�$���������]� ���-��O�ݑ�v���<�x���P�s����3B(���_�n�J�ߠ�5D�cQ�t�K�1)��	�9�j��2��b/�1���!q��:��9��F:����a@����"�	�蝶�{��L�Ȗ_��/���Z~��� �>i���-�} �^3u���
΢ ��oKe!�T�00�vMjU�>_ԗBIM7�{z��h��X���G���襅���?(yQ��Ϗ.Wg��]騄�)N���AR�S���Pu����2W�p��kGo�[qn����G_z�����܈(r^�K���NX�������{�"�2�X�cz�E�6R(�@�b^��;���{���<�kt�c�UR�I�)���z�&�m5���$wL=T�/-Xt�/>/{�U����2���&wķs�x��Ն���i��(~�,���2�L��1^U߬��~�wx�˃�bܙ�3�+~(�z{Uw��*�UV�?�3�%ȸ���2�6KZ���݂�JY9��0��.�e�V
&xu�}FT�C���|H;���¾-�g[��yҲ�J
��/���g��M�7�l�k"υ]�|pʇ��~�}�b�O���?�hS Z���w�}�;��O(P��!�c3/0gٜ\��Nק}� ��9����t�덙��l��U�������WSTu��[�-�<:�Uy�ξO�w��ڨ/U�%��HӪ��ݥsJ�������Ss.��=�C�w��-��|�k�i�Ll�I���i��KPw�����V�L�7�Ҩ�l���{4�/j�x7�ރ�'�XObJh�7�(��&�A@����?Q����-�����n�N�/�������v���~ ob���:�/:d~(�ՄV�++��NxK�4M���*,c�CvlD@��/>Xo�A��t7<��q�=x����>�����M�����-���֌�+�z����Gf0�*$���D�k�6 ��q���o�`-�4�t]�M�!����$��x؃Z�J�?�����;U���~��w�j�/i�T\�F�p]���h�D�i�F����AS�
����
Yh��K>� #�O+iZ��<hYJݛ�Qx_���mߎ�X-n�%�\�X�N(
�u�Fc��7����_��F@���_=q���S*���r �%��ǌ�P�Gx��IM��4ˮ^�4ؖz�6M+C���_=\ژA�i�>e|����+)����SO�n!��1�:-�/�ѹ�7������{�3_�|�0!\S���dI��=>)q�_��Vx$��[�Y�Ϋ:� ��;�[�Χ����t,F�A͔����8��iy ���t��f;]LTLSQ��j@-̿*��	�L�D�B��^_��/� M�����)�s��s�I��ۊ��
����27��\��6�":vV7||;��+U�W�)����W�����x�r(������d֧a��b�+:M���ճ���BߕLZ�E�~g���i�5rT1�����v�����'��v$>�!���$��t��Vqm�;|e�x�x� �K[���8�wlM+v�]���'���Ӯ^v7~�?׿f�ܟ'e7"&���	ȷ����BX��_������_`ΐih��D�YDp/��`���Ŀ�7ȨR�Iս�=��mӛ���Tay�0��j=jT�5�`�~c�;s������&�j�p��圃�mpP�M��T׻>>�����B[1�o��%՞p/��ji��y�׫�ZH�(Z����
\�6F%�ۨ%��H��$ 'Q�ϣ��;F�dM=��9����9��Fhf1�r�a����V�(�l�u)��a��`����@uХ�u�`$rf�Q�^����=��U���� nB;N�N� KH�e��6[��TA���]1�$\�.���w��.�|�[J�1dq�ZG��œ�i�e("��'f�R\b��6���G���~�/g7�JɌ��P�z�[s|�*��g�P%9�s �3RM��7$m�'�- ��U~D_� ��w���|�k �#/���5
�������*(�{�Q��`V�#S���'q"��ѵ�Eg9������6<�����2�����l���b3�#���E��p�s��ڶT�m�mS�:=O��"���82k���]`?푣Yq���q�W{�?U��a:�?-W_�wN��繮���խ��|N+�}�,�����LyʟՓ4m.
Z94��-z�ݞ�55��a� <�;a���s)"s���MsX܏��p��P{L�Ju9+��Np�p���#6(ab�����=���?�t"�I�R@OΒ?S��1"#���tT��)N���b��Ra8���,Ò��kL�� ;�^��b��e;����}̣Oxl�"�Y���K�7��y��+	_�]7��?*������H�]�'��S���e�:���%{�4��fwOD2}<md�)$8�D�b��TT^��4��S�w�o��D��V�;m^J�{���m��97A:�����,�/ۑm��2�2���Fy��i���X��N�޼��yo��-����g\�[��N�գ�R���r����Q<��r���0�+o����[*�¿��t$9D��S�:�DB�:!��;��<�h@�=i���YӗM�����Ea��Z�-�
���������R��4�����M���~�~ܛGE�8`��xL�?T��ez�l+즫c���c�TG^|����q
*OF$�/� T���ht�d�-�\��ίH�f9�88|#S�����
�+gs��y{q,p?�\�)EZЇ�u��T+�U��f��ek	�گ���<=��,9ر��.'��Q@�����n';4T�S9$��9zu���.l;�r�@��z�~_oS�Z}I��K(%gƻgz_�)h�'=d1�1��n �j�k�3�>�~L� �S�?��P�^lY^h�I"h�$!�B���^-.�c���u���x�J�@P��2[�(4���O2*_����y�8��� �`	E��b�Fd�uofq�\�]��R�7<�`!y�W�IV喏�c�=Vk��vJP�J�3X1�ft�?��{{�䟘,���i�|����|I�x
 �}�G�|y�D��us��q��0*?k�9ۜ�(?#��\�/h������jN�NSp���s綃�ʛ- ��j�tbʈ�Z)	�?�nlKd_�(K� ���b�D�k>�L�7��r4�^>�PC�4�{���$縎|���˓Lr䇆	�D�O�}�>���}��Wѷ���s'x��L�਌���a��I���}/9�?���w�~�Zw�1��Ѻ�r�?�E�E���;�Շ������L��Xw���'�;�_����Jn��Bf��a7(e��]�`ա%3X>�5ޔ�mY3�X��A)����Qk�EF:�����ڢ���CvJI��~����<�(I���ê�._c��)E��Pѯ�
ߤb�2�[�B�9j4q�I^c��"�:�s��@ca���i�Z'ޏaHMI+Si��}��?N#ܹ�L�a�_r�.`���gVB32�>��@ךc�!�S� %ebd��ă%NX2�����aa�	�.���ݵ��Nw<YUꦈI�F��y�}T���cLD;s��A��8�/�1��?6�?�b��3,�f�~�K��������a������A�i�S�0�������w��mwP]Kg����}����TYD��G����Ff���e����M{����� 1f�ެ���v�� �{䅙�4iA�AE�ϫ���n�į1� �K��[��KHD���N�1���V���� [�b%(g!����|��^�S����^x�g�}+�r�� ���.�&z��J1�ػ�-1���#q�#���(���+/�%�]I����h�,Rx�J�4�(F�f�|�P�Sj�s�g��n���0����$�!��
	^���S@fl�[�Ǫ;Ѧ.�\�([r<9������w���WT��r�~�|�����*�`�wz+F�!���M�4C34��q3���;�{t� �n�U�qE�!\�����XI픠R7*���(4޵���#��/>>��b>T%�O�N��F���yBE ���;�̐YS���������n<P�eCLB�ɷ���{��:qzvb�h��/�ַ��i1�N\�?�mN��RVJ��#���b�YJH��P����!��ۢO��0�U���/�,�}���(��@"[.��{@�S9�+ك��OhL(�L��ȳ�D���h����Y '���zN{�;�f]�?������MxU1�$�T9&H:�A�(*�S��]^a~��
	�\������E��ri��a7a��\�����_V=+�◃J�`0S-"f���2D����7c�n��ؘ-c��m`� .���a�R��	jf���v3��H^�&e��v�F�
�ے1�ݽД�����-�Hqi{'X��ᮙH�A��O�i����F7���*�i;h�a�����ڞ>�=�5#��7p���s�Q��y�(J�Ű�ϘD/���]!��Ca��@�z�� Is����C�����S��
}fE��z:r�1��/�cP�n�5���
ob�������M?�>��N�>�vĩ�6�����&*Cal&R��x�f�F�])EIYȇ�%��ʷ���.��D��n��f'�GB_�Wn�0n� B��y�P��~��|Գ�_��H���Y��[>���]�Ig�ԓ߃�����>��@�$�$��~�K���<���H�_���m����C��0�x��ۗKޕ��D ���L��ݯ0d�y~Mc,��f_z�ԩ�w�S�����t��_��3��Go��T���{�<"x��rq��B�����.x>΃wQǤ����%��|����E5 ?�7�c)�z-��)|�l1pG�{�;ZHX��!\�R¼Wq�b�<癫Ky��]�r�I��w�3gf��¿�����*�{�����{�d���kҭ���Ԗ�Dl�J�z�|x��/m=MTy�R�C����@�ߑ0��j��!��:�̕���n�[��Dx��]KT��'�t2�/�z{�7��t�[�#�23�yK�	���K��k�pc0���ߟ�{X3�K��c��߂pe~mj�\
ʸ����-�a<�=����ܙhH�6�N���XL<��K���oS�*9�6׶|&h}������w`��PY��e<�˨��P��H�*����t���kq�Ʊ���,�Ā:��@~ں;���J$�ٱ��(h�_!��[<5�O��O�FO�����*W�_#�P��u�q�����/�� �8*^?�|&(���Ye�-�1!����4�|�1��z4��9K����o��A���<>ؐ�|��!��o��\GiC�<��`8�:JSkԱء�0�ޥ2#��Q�*���Ug'F�/��J�<���u�#e�ƪq���=6�+�O��b���Y+�g������Kf�U�"�<�A�j2|)7>gd}�]е1��� ��$���2�����w�a^�9657�jk��6,���L�V��E���W����xpoC�`!��ӌ�}���&����T5?�Y���랕̢�A���N�&�m�#�L;��v����J)�m����	T ^�8��G�W}�X�m��)���L	^2�����YOȝ��Po�'��u�����u�F�V@c[�g}�g�n,	h��\<\��DL��en����M����^�O| ':�o�QnQ��ši@��}�iU�E�����P�!/G������%>���U[��ː��u,�p��!����fZԧ�~�1�)lu�e��L%���D�|�+Ƚoߣ��5$���3���-ݎ���aԊ���D\�r.v�%S�Ǉ����$mI��7�ư�{���C̳����?l1䵙V  |j�g[Z�BP�n���2w��dF�gq,6>�Wjk�m�K���7y��v t�	'�E?�c(��f�5�AP�*�k���5�Q�e�eDr�,��U�� �D�ݡ�ݫ��(U���������Y����֟�[&b��+��S��$��D�Q�ܵy��w��|u'.M������J{�����E�ox`z�<�M�:�1�&�}kf�������c:˰XP���P��I!�
TDx��2{��Gn�vs-���BG�����؉4���Go��j���>���2��0Q�r���\��|>���[��tϋ%xs���l�"��{l$��,]�lt`a��8R��iedY�g�����R��������b�%���_JZ#3���o���lY�(i�`
�Z~�Ȯٙ%�qK�V�V[�N�,q{^ۼ�6/i�Z�Ӟa���#x�J�v�ln��W{��l��S� �:	mۧ�e��W��X�Ќ�,~��+�^�/>�a��aR5|�%��z��޳,b��~H�v��B?xj�ۚn������Q܎�`�/��z]���r�Y{���VH����0
��'�3nD}���[q.*J\����J��Ǌ��V'���1/]5���|����4�ӹ3M���!��}�L^-J �N��9�m�x���!\<8���˜��1�:�c��b��W���(��c�5��@��Z��!��)0@�_�؆�)�x�_��r)}5�q����c=��n[t߃����Ě-��g�?�)|�I&t�⨊.k3�:���#=``M4��iOP����̃m���D�ǄJ3l���)�LWqvR��5���'�IK��� ).,�^���YYbv����@��=p~J"{T *�Ӄ�N牱��kN�Wo1[��(��;�T��&�r���@���t�ѯT�?�K�N@z��)*�z���e)Ջ�B	�h� ��_��D�ʥul]_��X�v�F�u����6XLnĝ������2N��p`���Ԛֳ�#��!Wnv���p�Usk�\c�	��Js}�/6$`gNk��A+a����~���������w����{���YxT	 ���Dy���(�m@�k��(tͧ���b���@��%�{"gF��a�]���=�"O��,�k���o�W�b�`�G���j�&G�'F� (s�� �O3��H�\�=���#A��qJL�c���l��m� nUnwt���ӽ�Smt�׌���i">X�z���8�9wb�l���h�Y���W/���IF`q�{��P�;
�ɶ��w��U�����$�P�����+��~��iIa4") H�)J(�JI��iA�]J(�ݒ2J�a #d���3�������'��������n��yd�a��vc.Ӌ]#6Ǳ�Ǫ#�f����_U�6 �ᙔV�@H�(��*Ho|L�� ��ff��C�]�3��A�&FE=2���}��%���Q���"ERp-�V���V��ڽ>��1�H�����t��ğ	I�۲�	�`�QE��X�vl�ɜY��ڨ>�m�,���
H�k�>و�$���F��Mb��cxQ��-;s���A03� 38�0'�i�)��	/ ��}JTԏ8�{B��O�a?��=�tJɳN�����6DR� x�q���f	��@����鷋� �m�>��& z��&���r��t���4������/gg����ʏO��qLS �?��2�"�<tRP��\q�n�ǌ_�4�IH˾��􇡞֌8 ��Lc4h�
D�Q �X9J|���3��"�/~А|��g|��O^���w�bp�&�V嶭f�5J�Rr��y���q��S{��兠���tBE+,F^R�[���-Jc�eo�ar��
vn$�y�����o{�`G�����8vA���>��w.w�X�`K>��r&�rM8�n�m��+�^(c�WO��޾�-)�����S����_�9�4�N�u���e"���?9���2�H����x8(��Kŋ��������7`n�c�+j����J�(��r�X�t����N�>��[����3�Oe�����p����,��z;jw7"��A���@���m�T98D�.��k���F9�0F�J��ST*a�%R�V�/k*"�D�����F�&v$A��o�Pox1GӾ-�c���mb�65��F�fP㡞8���kqA�~�&��x�Y�	�����u0<���#�ͥ�Q���e�w�-(�u��AK=,ܭ�m�;X��墖��s�W���2��k����HSe��%ҭ��WFR������֤��R7�c��������g͟a�:�T E��ϴ�|��� �&��)��$�e:�	Zk1�{�����`^�b2s>���N�v����Pv� >*P�eP/�pp����
I�Ύ����� ��\
�#�/��Þ�o����)֢�݆R�Nr��'�ucOr�P��}��T�聺eFdCK��g��K È�:A�>����S�B#a4?���jhl���	6p~І�Fh��
��om6�DDE��:�h��=3*�3��>}Ck .68�$Q$?�;J\?�����KQ�d��dܦ�CL���Vn���+۪dJE��A&� Dɶ�Jq�}䎧��lӇRQ�\�(������L�{K���&���)nh�'*�p�Hg����7 -e��Ӱ�� �=���~�t���"e��Ŷ���~<X�jI.�C�����k8�L'�Z�%�I����La�����̡ߨU?�}'��P�l!'p��%�{2��3TJ \3Z"s�./�<��t�������D鯋 *7Z\J�<lJ����T� ��^�SOg�9N�寙_�
8YMH���kI�J4 d�����ƪW��zp
:W��4� ]\�(`1���u��  �1���7����b�������,T=ݢ��n�Z�����C�5P�"f�	�axлLʐ����Sy��NLP�L��F G��rF�@\�[�"R���NDwU�./M}�m4(%}a&* ��nc��]V�6s@�JT��~��9c%�a��5��� �$���pN����������3�I)i?{�Ԧ/����q�M�hz�}��MU=bJ6wT��pa�x�z j�G���A�Y�}С���8��{(N�� ����vh[�Z^���8A�3I<,WB��$��ћM�!��>;)Cqy#���F�8F��Ń�p9S	�ѧ����/�f�$-�Y!���v"�C���̀()KVy/��6���O�L>�2i5�<�Lyy�s=v�� G7���UW��ȰB45u��k,JtF@�� :���G/�@H����	�\WUؠ`��5^��uشpsK�&�����ɔ�B 	v,���M'umIء1�]�'O?�e�I:���EU�_`T�6�������9�^�i��U��f�L�ԯ-R(<�o. f�v�3�����9��KG��4��/|*��P/2���������9� �T$�Hq�K#w\����b�:���n8_�]{nUY�Z﭅1�1�$a�����ʁ�J�S�Q�g.|W�B��W"8@�n�u��v��<̈́���B})�B������]"�R�qA#o�@���:��9�xə��o��y�[���oQ'��燀\���|7���A�N6�*�[Cdΰ�b�������]��_��9KͿ�jO�8��	�O�_��e�uco+J���fJ=�gy<������b���l��B)�����I�_�A�E�.S�G[���>�Nc�xԌo��M�2֏�����:qo�=ɔ�l���[2���&��|t>�ԡ���Q���h�t�-�n^,�(��	0��T�,�����B�S�Kv��x��N����&<u���cU+�~W�*��V=@�N�;�1��S;��j\`Bi�U/�|d�|�l�5R�����z��0��ێ�n@�4��g�85�N�8 ��O�N�u��W� (y�W��O�o�n�%���0+pq佉�^:F0����ʊ�*�J�O��㺫�Z�t���4�;�l���ѓZN�f����5�����k�ɬ]��v�_�L+��v�ܺ���_�_������%�O3i$��@N�?�h���Y��<�q1��ԑ�"��g�HEO�LԽ�e�ٮaj;����I �&F�{�J���E��M2f��RR�Q�.�P��9+��q�ϭe���)E������R=���������b����p\͔�wz�]M"��[(�i���Q�]~�?���iw����J����7lda��!d{�^V����l9�6Z�EK7��'��B( 6r��]�����s���*�N�?�a���[�ɺ���)%N��[G��|B�=L;��.�/�Ё¶�~5�
��(o8��[h9�EM~����l�s��Zu/��6*�C�����0���Y��c�K���뻟oUǜЀb�$|��D�)�r�y�c�1\h����JP'f�����N�lBƸ�@ǔ�����(���с.:$KvD��P\.HX���.�^�ɤ�<Ղa^a��w�V�}��LW�5R���a3������K�w��s@(�Cg�2���#�'T��ޞ�8F8}������s�%g�<��"�ߡo��x�s8��O�4���;��X��A
`�qu�D�:���'��Ȯؠ�>�Ә�	���
�fL\��=�kpK.�@)�Њ%�_gCZ&��L�~�`a�
9A7��DsX��a[Xc�����r�1�}�u�K��)�g�f�>6�4xzBu�w��'hs��g���V�*���%�n�Mb����������M��g;.��ft�%�z���d	p����8�܉|/�`���Ʋ7ځL���=��<��b��单��_:���c=#�?�T��	�/�K���OŃ��j�[�?���Ŝ�ZA��^c�'H����������'[\�T.Ee�k5�C���������b�3�����=V`����o�aٌa�fm�Z���Jy�s�|d)�S�(�Z���nY]��EN����,"1�œ�صd��9�j��}�/D�o>�Pa�h��R+8���%��B�y��X����&@0i�q)R��R�1U`���\�6�����Ğ���t��?H���L�!�矍�g�s�T)��%�X��~��ikU~Q�����\k����*x�K �o%Ћ�ć�<S� �^7�̣����?�>݈\������Cj�Z���7Y7��75��!��T�����\��=�]O�*)@b������9���d��P�F�F�/�'<�d0��V�,o�R� ���lυ�i�����ɔURV��yFL*���U���|c��>$2��Q�#v�_���I�L��[�l���d���M6W��Mp�M�Iu���q�S�}���nu�O �f&4�k�J��5��r$cVȨ�-��e�%��G��ݗ�	㖆��N�v�!*�27�<I`��VO�d_�-LG���/!9i�Ć�ߥ�
��ϫ�-L]�`b���3"I�u/���A���o��'P��{vJ]�o *��ۜ��˯��4wk�t���FUnl�dX�(B�2.Ԑ��S�}J���n�w9���M���:!�P�$��Z��ư�J���5����I�����oǍ�hƺ|ȼ�0�>B�U�#�8�ԥ|l�!�Q�`{�Yyas��'�J*�_Y����)Ǥ�H�W輸�߅��`��3��&�A��n�	�0����9$zԱgi�t@?2��҅����Bg�dV"ZB����lp�=�1 ��1��܌���L��x��*�Q�"Ն@��Н2�*�f��7*GR�M�}��H����x����d���~��fc���W����OCVjO(��k��g�ߗ��f�#xp���;�%UNc��{#�Ipڈ�%	А} ��3�����q������kD�����̆M������RS�*�8ރ�~��g�W�@ޏrcy��۲n	ah�{D]Yx�]{���i!J�+;�3�}���\ɱ/-Mf0��I���%�����`C`Q�V{�E�����c�Z7�UC� �W��Dԗ�hb�#
~�b]�4�E������11�J�i;�4��0�Bj����嗻ڱWW��R�j��4'�h8�ۂ��:�i��D�d=>*��1�)�6�|�!�v�s��z��t��ɖ�u��N^��g�O��D	D��,�Rw���ݜ�g>�Pr�Q7��O�����21�'x�Z �UD��7�4g0o9��$����-rAc�aT�`U��;�5Ÿc�^`=	t��y��+�ٟl��4���E"����.`�i�����Y&��c0.u9��Ī�����=
������N*�z��a��|��c_8���FYY���r��㊬0�߷=���?zK �BaX�G�!�,?���$��p�jO.��9�fA���
�y}�b�Ϳ?|BU#�ϣ�fE�[.�
�	��	�.�y��b��d��&T.�D/�<�'P�{n�k� ��E�zc�=-m��ܼ�u�:O��.%c�q$Å��0����f�����%��4��;�����S��LQH'��h1�P7v�Z-�[���ij�/oӣv���Y� �*���B��<�%��B<�y����V��p$E�k���{jg�.���Z;Ѽ���>�
����e�w�RjÅ�E���ƹ��V|��0b0��J[xc$���x��i'hR��G�~po�h����� ����-�2��;���?.�Y�����9�������.��H9Y�
-��r���i��R��^�0�%������~JP:��{��@����:���A�;5}���&�g���,	s"w2*D�Gz����� ���jÏ!��Oj�`X��j����1̸y�������S�����!�B��Clp��1*J�o#�8:��4$��q��K�ŸX�qaw�5��`P�&�B����L���OF���?8[����1�>_m�ݵUV�z@J��� ���*?�3ds�}�����(�ҳUVU�;	�H�!|'�����f�"�v���7R��\�����J\��j�дx��x��Q�1�����T�$p4��FB�3��PV���m)x��3s�ķZ�����='ӂ]e���@���V�L�\�4e2�x_�!��d��і�2
�⾬@r��j˙s��o��R#U�5��W��`" Ł(L41<SZ\+bh���2�[! ��C�(Vϗ.�G&\�	#�[��!	#CqJ�:��o�AR�zH�Z+�J�҆%b��ʔ܏�}G�!��*�W������������y���?â;>tI�$,7^��$H��pZqF�=2�7�UU;�Q2�"� 3U�C@���G��ՕY�q �����c���S�Ԉӏj��}�Hw�^fg�Vb<or�F�͘����t^~���J��_�}���_.#�Oe�K���Ҽ�B �*��t�K;��G=/t�\�7��ֲk��QV����r��kL�Zт��eqn{5W�D��S *Fq��Y���)�͚������:��L��.GF�/ɧqU]�Dh�sд��|[��@����B���Zd�w\�@�����o�5�	�x	>5�F|��M��g�	�v���6��!�b���k	��	���O���o������� 4�j�ϭ����ʸu��#�mTWT�>ǩ��X�8�p#�S��d
?���Z�l�kJfx��"M2����ir_�%9ȇ$wӻz�#�;$t���������ً+�t���BJw�0qP\�-	���C�]�
�
�T2�y~U�.[--�}���\�LwYn���8t�3��xc����l:;4��'�5��� ߦ���V�N�;�V=�=J's~h�� ��@T��2ow�/��`��8�³�\���SU���'�q�#>|�гn�NE>2�i�4�����3JF�y�dw��L�T���%���˿�T�bU�Ϡ����ҥ`��%2}�I��R)g`pX�-�@-�iY���(5��2���@#]�W�|es����g��Π�A1��X۞���%H�u'�yA�ށ�`/��xG�Oo���:�Z�zy�TJ�9(��rS���;���*�Z���.3w\K�Z�=#M�؍y�h1C�p���ˋ�kMx[��G>FDjF�5�����S%u��șV��\�*/�v.]���q}���>�ן *v��{�@a�o�Y�_��Х��+���z���%��p{��.P됴ά$�N����]�D̮��JU��
���ؒI��/[�(,�92:����12
�ӣt{ӘhA `������|�G�j��<�:?�dF
{Έ���L��Z��Ξ�;�g��
��#��ɜo�e��z3&��j�0�i��CV%�#:�Q%��<"��� z`/�c����%�w��{�Q$w�.ð:�
=z�/�����q�@acwp���k��.4���*5Ӆ#r�!X~Q�"�{�Hb�!������@���g�����vm;����p�a�u����$��_#�B|`��%���IGza9��wl@�Oa�o�)6~&�~��K �U���ᩙ�:��H�{S���NFG��C��#�ty��k��Ʈ'>��[_U�_��}��3��.Ξ�a�W����O���7�,�~�]º���;�W�JTx@8��t%�Y��z���ms���'�G5&,k�IF�P7���s��νU.��t�S��y�8�]�/�eP�B̟/Latk۳�5wP���,���E���N���kouI�����h9v��i�]�  Դ��g�:�Bk�;"u�ŚT]�b���/�a���%�R�o4?�#�1߅]w��g�Ef46�]ât��4��7,,��z�$z�Of+]��=�+jm�7OTw!sNF�j@�b�#W���b���Sk���]�;*}m��4�D����/V.${��lI[�A��3d��-��M+Qo�޹>w���B8��FY8�y��,eΉ���yѕ�aاՊB7 7Knhf�h�diڮqp*B�˫?K�u��4��\�{�sH�h��(n��d�W����{;d���#���W���Ş�7��61��EQ�2ׇ^t�{S��+��@��,���H��B*L������t��X�S���1}������̥���tS!���2[��A���Q�QO��P�N�u[dJ��~�k��y����c�H���)�G�8$z@Ǽ��ie�ݐ�ɳq�[>3-��&:dT�*GkE�kMݥ���-��hPHMB���)X_�4{�ܯ4��J��,&g�@���v� ���i��%2���AJ��b$�}|u���-�L�GL�)Y�?X[�����������߳�;�x��)j�œ�۾)�޻�U�{�t7<�:jٹ�]�_���
G��u9�%\���P��J�B��u'	���'��s���fHJ��E}�!�P�ٳ�dn�҄�[x�E<Х*�iq]�|PU��Q��a�$��-�ٚٽ���VKa�� �\'��i1��>�H�Ի�%BjǦs	��3��
z��꫃F"���9���S ���s Ӆ��2��<��\�� s9s� [?�AM��Bm����:ّ�3SEee��D[������ج���'�����"���!q��SQz�����Bw7�j��r����k!�ōcT��.��|��������l;�6F�ĭ�(��KdJH����߇s�G�m����ieFk�U���nЫڡ$�Q�)�S
�����;ǲP~_����dK�y�Ui��s��:o�����GA�U�ݝF������GDХ������ �qsN2ta�v����~��F뛑��	��o���.r�+����!�9[�:�N������o�o�����'��r�M;K��{)&��rc�2�'���M.`.��9�AѐD���������%y<��c����9[����@��C�K犚MGk����QIA���������~0�Sq��6o�}3z����[�/�l�v�2K�@������<|�/�kh8��fX�P �U �K��=�K���G��77ݳ&�JA�p�	9���Y�U�I���T6��	+@�a W����CtM��#y����V���RT���UY�HU�}���p�� �bp?3���:ډt�`��7�Z���=%��7�O_��l4�|.V��{���^��¯![��{��9���:b�Q��b䜃ː?3q���j�����B���G_]y�a`Wv����y6��e��l-��?ev��8��ds��2��q�lP���1JB?�u�&3�.���Zj���T`��U�3�ր��w=�, �?+��h�ޠ ���Tgf-���Zr�
S�~���>�h���>q����j��Α�E|Hw�ȁ{��T�r�g{�Ƚ�sV��_�ʟЛ�/�p�7rN�=�ۿm.pW���-%�]x�W�9�W�S�T�iГ��\V���� s�>�}�tպs�$��͸=�&�G�q��ȝl�x���`����ŋ�����ܶ��8���fj�4� �ꢻ�(jO�
����.[#�[{�	~�t��{e<5w����	�X����o�^f��8(�e�;�Y�#��ɡ�k���7^�9�)]x�9�^�cB���8�iY�6G^bbzVW�F|�X�>�g�b��zĞy��j̷��d��:5fCL��x�C���G����yKInHzg�	����h��>Ru�q�w~�Ʌ����j47�}��0�ͻKNȜ�y��2V��Z��5��~�q2z�a�s�a�`��v�p�[g����-F���';�����.c"$��g���ãV���h�3#�m�;�#�ɂ/&����8����O�Qۨ3�⊛O�/�KpP����g> �@�2�XS�,���^���e�l��K��/��!��_�RO��ܞ����!V����,\��Gq�bd�-����̲��9�ǆ5_D}>����^�*w�,�y�������3��&䫙4q�C�(�ΩK�U����ND�E�s8Vn�����B����gK?�����	���F�k
#�P�_�=��:t�t��|��p�ԁ�-�.�Dˋ��:�[�ǁ�TFuQ���F�I��y�f̙s���Ĝ�U�z��X���sY�������� �(����QsyQ��bD����ȧdDξ�uBR.�<~���3��:[M-�/]q�f2��K��<��/�eZ>v�h�l�߭
^U7�p�+�����K�ώ��1�uC����k�}�\�Y@�ޙ�
"� 0>�dΨd�E.<�� �����R��n7��޺3�3�(��O�o=�����@���D��n]Dܝ���pu��#vN1{Z;���!��]��@�����ʜ�px3ѹ>��ʐ��l5�~�'��VT��M�6��HY��#��|�Sl6�*S��o�UmU���-58����c@���a�"W����W��Rl���{���%�>�U�[nAqtae��ˑ�Z��	DՕ]��Ƌe�O�Kg���%�]���lO������`�ݟY��N�}e��~��i�ڸ�Ϛ_hޜ߀�N�'�l9�+�@��\w@V�.y ��V�$D)�ۗ�!��x�#j>�@.����2;�_�w�88�o�훪$5~R�u>�T�Yݚ�@�� {�M��=���e�<���7g&8��}�)
���2�Q�`.�eჾs�Ф��D6�5��lY�Tb��'���L']=ؽ :x�
���큅<�re'�K�[�֘��o��A�t/zu�_$��L[��=���(��V4ݲ����G��Au[��Y��� ��d�1,3"�x�$�`�"<(�U,1ڂ)�H�N@���r�;�Ʋ�߽ ��@czT��2C@�%��5@�ز��Mj��c�(���߸����|���x��]�l"nh�z��z�go���iΥ�v�j��l��"ۈA�������L�j��h�J�Y�y';,:#���-�i���g���,Jo��-?�*�l�:w龲�
��
���j#<�)ظ<��Qf.\<���
�V���~g�����g�k�`�b�e/�������{u��Q	��Vy�v&���]�����e+�7�B�<����ۧ7�0�y$�[R��A�������o���@6�n�|�g�s��V,`K,W륥G���8�}�$�	B�ȰLs�YVu���ѣ�㣅6:�z=���/�xm�gA��*C }�ZGԕ�w�X"��;��v��5�h���]�/�9w2�i�Ơ���kG2?@¸�� �#�@�l4�ڀ�yۋ��4�95������� |��7�֗�_���	ӛ"rr?��8�fS��>�d��>����/CcZe����	��c�&+5E��<�_<.�L㣱�Lq/ �x���?��9a��O�)�i
k7�f-��\	�mG��^�&��>���
��&z�/B��>�Ӓ���9${{���6��Nd{�2�L�?{��K1yT��,��f���D���?�V�s��e���c���F�<���	��w=���2�D#7]����8�+�3-��'���o=�Ix��s$3O3Qe�A���i�]�u�=߈Q�2r��]ժ�w��:ՙ�u���3��4���D�i�>��@�r��+�~*���=dG'���/�w�7��f��G��S��iw�4��f�H��۹��<>�Xn�H��8�7Z��jr[C��G*=�L��񔦬���dq_�-)�I{���fZ��*�~��DUR�����x��ijt�l�6K��շy-<��G01a"��ǈvF���
b�
92�,�d��7O�OUi5x^e���a�['�_���F�Yr�V�,�tmǮ+P����z��U��|`ܜk��bձ�#YP�qv���T��="<����<�L�&�)ܹ��|]�~�{�Tj��۽9A*��ppfq�M��BN�����FT��ӆfv��|�B�Z�[K����� ZB���&���/��u�SR��.�	�X��I�-��o&O'�wc�j�}����B�l��ؑ�� ��4�X9er����suP6��raa�^�V�k���
\�z�(���ń4�iAjmc�{^��31��v�Yo��׾,�4f귅���炟曱\�:�,l���|��Bh���]+0-�?�%���̻�䠁?	���<��w/ �2`�Rm~�9m�*Y������
��τ��3��z�\�&�Nu��dIG��N�����[�4�y���{�xlH�ܞ����t?3L65�ڸ���<�hS����8%e+��l��E��%���1;?�ZP{@)����y���/�5��n�j�Uc�$zțm׳?�t�ϭ���sO�����7u�wRϬЃt�@
�10m�~}�����JM��w�ت	f�B��J�����	���M��9����@��@?y֊������T�{Iv�����Mɳ�@�{BxS��R�\a^�/��G]X�ݖ`3�N��Y`$���f\�^�:�A�v١����E�'x-ݫ�s	�mu�9�U������o��ԨIL�b�eo�r	AIy_}��==vJ�t'�<��	�lгq���fo:+S�KW%�%�1U�0`���P�*����V����D���j�u�,%�i��$UI���0��e٧{~8}�9 �����gH�r�={�U��r4���MKGSbՇ�`���$��x�;���	��e{5(�*f�o6
�n_E}��{����;�2Z��FNh��1bo;5q��G�j�kx�b(XcLU����`ʢ}�)?�H�1V��s`E�0gj���S��ͥ�z��9/�:E�f.v���̶Εa�����'9��'"{���D�Ȭ�(��>�R�*�l(������`zT��(,�]��{�BC����O~i�����a����seM��V��_�0�y���['�|y��s&o2A�?��OȳʷqmoҐ�@�Z`�Iنj����
$bbz�[�t�6V$���E�e��>M
zq���Qw2U�����y���M#9"�y�|��|vp�X�!H�?W�#Fp����)�Z`|ۣ��?���2�9%�-m~s��!����7�ۇ����<�[�eGUf6��3��T�k=�zu�aϚ�ކ.�'�"F�� �MBИb`g]��	Q�+���s�p]�!$Jp=�IĮ��0`[C���fB��&Y�DZL/�lXQ�`�)��k;�O	��Zg�'��[�\�Z�����љ_�:n���}��'P�iwnxiF�����S�GW���h�`Z��Q�\|�6�'�uf��K.e�ȗ�������:���c��o�>�%�h�X�����1�~c�]N����Hƍ�S_s��'��Mc�89A�|c�2���o1������N�r	Hi~[a&UN`�P�	{���⛉bH^~ף{8n�����o,�6_^H�r(�����_	eV�ݏ�9�M�t�aY�l�1B*k[�`5^��*z�A�,ާ� }g֍�a}��Y� Ԍ��j��T�Bn�*��܊(�<����R�����d ]$�'{�c�������N�X�_��
o���ȭ���%$sXn�&����Y��̒yg1�b �~���G��cj���X+&�`����O�=Q��_+V4�2�S���|J��_�,T���<y��ςM���?'v33��յ�(��ֲ��RM�ʧ!� \����Ҹ`L��������/�V�Oܚ��2�TMk�؎�*>�r��'j����M����4�؟�?iZ��y(�J�>�3K�� KR�,�-�3q�@�ln���yD�'4�Z2߭F�u����7��6h�g^{�@7c�9*@M�.!?����Y�R���<�����>WE�o�l��vY�X�C��X
�����V���>�H~�^���k��.4��֫!3Z�{ɁH�*K�����۱�sNg������1�qѿ�
e?����V����w�?}��!v�+�2{ 0�s��S����w�����b��^�q���)��ݬ%�(b�����e0�r���2,�����jG�M�4U]/�qC#�}#{��(�M/*x�r/`���?I.4�}�j����R8��O����?V�Ey�I��.�Fw�����,!��������c��I��)mED��5߯���� ��*{י	�vn�!#���(;��_��B���T����'�I<��}'&�T�L@1��\L��Q)k���]���@J�J���q[�9� j����&y�y���⎩^�f��v��_p)�t'�nF��#��V�l`C�W�_w[t�����g����R�����t/��c�@���� ��JI	�w�
�O@K��tZ�s���NMّ����4��[�q��t+	��fh��ٙe5�>׌VU������rY}������̓�FO(�Z�b^���_�� �cw1_	�L����k��1VES�E��(�m�>����T2�)��3ڏ+�
F�3�z1
7h��<�l߼|wq���W�{ܽ��^</Mf�i���q�x�H��$gF�z嫅J倹��X�~�a��/n�_	_��?c��&��R	m�BS�]ZQ��g�#.�Rܜ�D@�M��doo� ��i��r�t�1	W_C���LEl�<>�uH����q
���i����މ��+�gr�Vwh�^��=�E1������7a���-���v)}�"��ؖ��	���1�cR	o���j+���0�s�a���ܨ�k�/QN��\����.�@��@C��a�ѻ�S�?&���y����\f
Ul?X07��v�����;�-��Z<��.;o[ki&,�1�ao�q$����{4l����/bv��sF�׏�6���ƶ���n0�MT"���]S�$	� �s)�.��$��z���Tg)$i�M:\x��A���l����鵌`�뢫���U�O�l�O޽M7(��0xrqJ��\��.=�7�������gqt�=6�;7��\���P�z�C�+13�^��7�?�ҐD>�ڏx�o����w�6=v2��j|�>�z��d���@*��}�Z���駛9E�B���<�T|�t���>}�Z�T��F(���}R&P�p�1x��뭚�+�1F��t`�/��o��0����廸�������NQ�7t,=�Gc�9/G#9��96^����ɠabgȍ����L8�ã�Y�^�H�oeG#r�:�74"8^87�{e���ͧ_ߑ��?P��L�I����#�|?ԕU��ׯ�wB���Zn�ӗ��Woh=
R���y�4�� 7�� 1w�kE�5̏�п�z�O�ۿ��ޮ� �`-V"
�C��)J��ۨfU'��]qp���s~Ks3�ߓ�����������2]Y2�7MZ�y�׶������{p��s8�mY�G��hZ�u9������ѩ�_��ʱ�u~Ջ��;��� �.LԚ�T�,<�8�-����{��=��Ahc�C!}AV��`�^��M��bR}��xN�����H�d��<1�K���bORD�3'�bv�8y��Y�1FO<�';;L'2Ks��S���������x���W��T�kE�.�ƨF=��XݥyTɉq&[U�d�3"bmc��9%!�e�{�Xoe*���37�g%3!;�����"Y��6nv1�tS�tR�S`�S��HKQW��n��H9@��W��H��!�t��)N���v9�r��f۬`ߩ�ةbw��W��Q��}�њʨZ wwQ���x�hW���;D���>���X��#�"2�S�~z�3-n��ep/��8k���p�b������J]6��v���*]"{WR���#,,��Ȥ2y�6�X3�g��kA_>Ȕ�	��˓��H���$x`�@")?��R8��_)o��r���t=����E+��W��6�]vj�/a�v*]�t�	��×?�i���l�
�t���MF�'�|�*LT@C�-y2���W������T�T�>;~�����V�ߤ!��9���$�~����o
�[�L����n\���M�9�W�J,����%h�?�&�*&����s�f'	��%F��=,�v�����v$��J2�Ay�׮�4��$��$��슴5�$/}� 7��72"��T��n�{�=JMm��ָ�Bz�d��%�z�u�pfN|�����C�S��~��>�� ʨ\8J�]��]*�"7B��iH�j��΅��|��9�\�E~E�.l
�U��ӋA�[���6�6��¶�%������z�>TPƍ�O��rg���4�����_��������0�0��g�~Z���Io�?c�ɋW^1j�W[��ZG�}��s����#�K�T ��/��-5���#����)��Χ�^����FG����'#&s�ӷ} d�K=f4�y�E��'5yXi�M)�t[]��ĺ^�dw��;m$�g���՞G.ޭ�W#�M+�XZ�r�{�j���ߛ�W�=r�8!y�^3�lywQ�D!�88�?�����Ʌ�[�a�]�������o���+O^ur��0�?`cv��\�n�>a���o��-v6A�U.̥�ӭ� �oD;���sI�EiwoPvV��o��}w�+�GG#��&��8��p�>2t�P���ZQg����^D�Q��"q�Ϧ�o?���Ayq{�O�l]�3Ojka�{�u7%���5EDi����t��zvR%�<J��
�ߩ�����7Jj�xI��{VtLn���dy��&������|��/�����(�E��(}������X���%RN��z������n�'�.b��WŌ7��s� hs�������i]w��3�apq����9�z�CԆ�ӧ�3UZhU<�Vťxx�[}�Ql���F�����S�=�VH���L%e������P~c�N���ո��0�C�f�8i�>@�"�B�[P�O�L���5�1��/ ~6 ��;��L0��v|�Q"�� QT��#Y�]t�ىD��Е\̽vZY����XS�k���޾�[+��4���6�`���3Y��W�<L���~˚��&����x#1�Zz�er�������	���g�8�9K�7u/�����g�)���.�mq&��������<Ÿu�?;N
�I"׽U����h�:������I��Hv���S⟔J.�&�P����Eq��N�]���e&c!��u�ܙ��ʣ���Z�iΜ����:�F!�9n��.�?��,W��'�*-��]U�÷��9�u����0��B��K��ˉN���r����9�h�a���ݽ"2�c�X4���n@3e����*k&��h��x�c��|B^�c�6���!V���{����� ��)���8	�L�99)�e�sv1���L��3��oA�(��]��>��ʊ�?�p��`�é��/��^`�G���K�b�?��̺�y����m��yY�k���>6�I��X�fv�[�I�&�0"��=�q*�;Y�`�k���/,7�� ��A��H��`$�k����[�E�}��("��4�t+�t-"m �H��ݠ ����-J���5���0��������/��9g���u�:4��o��7�����O�'t-�7�o5g�� B��?��71�G����g���B��֡ך߼�w��_*Í/yI/B:��2�"���C���-��F��T��Ӹ���	�8�#��v�ۢ�N�Z��ߺ|�
j"����5,�(,�D��"�w�j5�	�v#�|5�a�^k/@7�']a�i�˲��D#p������,������l*�q�����?��X�WWd��P�ʵ��m��X��cw��Y��'�8?��ɯ]R����"'BaT���l@���I��ρ�e�&Uw�$��铹 ����yY�"���������{�r�e���8ˣ���jT���걽0V��L�����c�u�ҴJ�:0�T��_��-%��F�g?�J��2���Yi�=��WW�Δ"���A�'SH��sғW��~��
n���{���R����m��K$��<��þ����������� �Д8�g�k ��]�oc=���p�*t�Ifc.��`}���͌=��GEF6@�B�=Ƕ����1�q��`�� wS/^��믃i��'���g��/�䎋|`q��xY.2>Ԓ���|�'#;��<
,$�����z�{��ֿ�b�G�-��1�t����n���o4�%�Uk��N���[��Y>%�fU�ާ++���4�������	�ⱐ���gyg�ٲE68�g}�p&qyQ��c�1����?~�n��},w������<��մ��4���7R��0���`G�_��+���_�ߒ:@W��ݒ]���7R�p�d9�sְ����3���ټ�I��oD�H��Uro���r"�~��韩��x��M�y6-a���n`-����z|PJa�]I���o�!L8������Y��.�ͷ��%�.y4Q�TW��y��4��J��ޣ�f�*�|=��ԧg$�]��ه�xơ��(U��i�� ��N���B����A̋��ў%u��"���I�	��Q�%H�~�
�k}B�U�Q@��ݕ�􃠂���9,�ts��(,Ih��R��~���iS	��������0.H3Gr�aQ+5��):$��l�҉h�%�㗃�]v$Q�	�Nk���oN�޳�Bw�MD���ط��֮��o�2E�]�� �n�r���j�(���5)~���Ss��Q��y�T�~�߶�I�o����7�����O: �7�ۏ�1&-��&z\�wD�d�>�4NwO%�ơ�i^Ctam��6�rnTW��R��7�u��,�m�x?nk=�W�? )x&�\�MK'�𲄒��=	΋{[�����$O�@U F(b���0�3��˞J��'k����hܱ�����/������&>���5��<�lE��i�ZTm�h�w�y�[��L��n>�A�w�S��v�j�kԌ�z�I<DY�
�m��mH{��p�)9N\�t见.b��}�(N	V��u&L�Z�W�j޻@�ٸ*��F��)��f�<d+������2����,o�-!k��G˪m������뎧Zu~ש�9��0.Ы�{��2��"'Ld!�(��a?�
��?C�����a�:����ё��dުRv�3��lI�^�v^��C4;{j�*�c��k'����.:)̯yU����V���p�8�Ⱥ��r�-��L���m.}��f��\g �U�րn�IjىHzU�'3>�'YȘ�S��xF�GH�罀l���l/�ݾ=<�͸#��0 vͤ��Qɝ@�W��H.R���")�~+fz��y���/3�i��n�Z�!OdӒ��e˥6ҍ�s���q���L��[�v!�Q����%�[��ItD����hQ(!�|t�����ދo�JDc%��{�T���o���(�eLg�[I��T�z�AzN�B1�+�C�u��L��9nl?Ƀ2Cۡ�5M�z����0.���=<$������;�D����׭q��5��ve[��"X �z�n�N��#c;(gZ(P�Y_9H6č��"S� ���zF��~����R�ʵ%|hl<c�|̢��#ƹK}ɤ7f�oj2���Q���^��zӽҖ�>Tc�ǯ��L#7�H��Dk0�2c�^2�+[������j{��b���C�c���F��)�e�I~_��A����+$���+
��Q�r���� ��ݎ����6q�b=�Ć�iKz%7�a{رz�5}S��u�ݨ/��x�UrA/̋<hG��;L��
���^6S���^�+����Ä0
���$�Y����	+p��i�~@��й�B�=̨�{]c�o:�ʌV[i��*b���)�r��D1�r]X�	9U�2�Pf3�e���ːd���n�P�4�{��沵�Rieb�?i�<g����S��(�r��ۦ�4e���o��pP�V�5M�"���-�����-KB]s,}��r�Gg*X�M2�E5)�����G,�*�����_�F��#8�[/�Ġ�E�N�w�v;N�t��>�H�Ug%�i�v��w}������H�u�S���"l�����������&��ds���X�<� ���qF�\��%7,��l�������WVp���*�e~Q�g��[�m��m]��&���	vn뼲a���A���摊����B?��r��v�^B�;2�)��F��dH��ژI��X�"V��FLqt�Z��ZĒ��T��_�S^�}V����Y�-!�1_f0=��WxU���J)���Mc�TTo����P�觱��<��hRE֗2QW�Z'�4c������6�G��g��CV�o�҃�)�m/X=M����q��!�
b�vN�m;��sd>J��C���	���=�?�^���oWSu���b(��s�JRR�)��2w����w�����sI�f˹A�wn��Y��G:^T�S�U��R{Y 8�w@d��ɽ<Tz��L�*+���������+��^�G��A�hFg��}%��KN�&�h8,�%nlF�wt(�3̀���{�t�Q�1r��4�n���_��	pD�����Գ<*{���	����Ý���gN{E>�LdŔN�J�T�3�Ԃ�.���Vj�BIV*p�O�q�?�<e�?�%���f'�`.���=w7��.�:k�n�~ZPr��<3N(Xѥ8�2!zbwJq�Ί�P�^VZ�h�i[V�q��+���*~���Q,g���)�Ƚ�_��`/x���Z|�cFIʏ����A��l��o��I�R���m�A�&@�p�?8��"��w�����ܿټ�e��Ni��y�c�`l6����t�G��d~�kD	�$�����z�d�ķ{�o����l_'�~,�Qn�R���o�_,�@�_�9��F��ӗ*�Mi��7�z�AҨP��]���?o@�IgO��]�~�W(���GB���x�1��4狣��Qsu;e��C�H����ϭ<$�]<��C��\���謸y�Pu˦�SӅ5����6���BW��Y ����@�e*
m}�u>���pZFEOQ���Q��4l�Y��K4h�E�t?�bɢR��g��sO�@-�_ܑ���o��C7��C��^�Dv�|J��%�����h�\G���6�f-�d h5�9�;1�M���/�1�R�|�_��$�ڤ��Ԁpi��ť�X1��?�+Q���_����,�����E>��zV�zEk�v)�c1�L��s�]�}��Q&-����\����1�sq��G:Na�H��$Q�#s��&f�(�t�K�,�^+X��Ԏco���g�Ijc"�갲X���
gs�b"w�y$._Z�e����R@p�59ަ�����������_���ٚ�8� ��X9ï�� iY�v{^���+Ò|sR���3;�
��Q}� �\
��K�l��9^8�E�T�W���p��j#vqj�����).���6$��Pao�P�Z����UQM��%�t���&��8�w�1G�r��v��ƳH��V��'����].��ҜzMT�MW,��VY|���;�<�F=��MPQ��e}h v��8����Mәo��s=8���Jo!����p֖"����?4���J��v=)x���a[�g]�W�m�<�G��2�nLU˜������z\PU�Ѽb<�\�,��#��`)d�x�L�]}��߭&���Z�j_8�*�]<���9��.��n$O��rnq%<;+>��5Ar}�/�d�%F�����1k��Xx�߫2պ{;4�RBR,���Uk-�[I\���r�T��	;г*�?y���W���ad�n���c�
������O�m7�Ǳ��ۗ+��u��v�Uh"� ~��Ī�29Z����[�������jXX��kJ��+S��Wm���wps�$4O�huy�d��A ���
N���Ef�'jXn�����Z��$6.����+�Ӷ{)z{����Rd��2�͍B�bMצ�w�m�r>XY���a�A؟I�7)�d(f�����b.�ͷ�5p��5R�m����1JdFQ��{8�1���#�W~����u ��0����ϒ� _C �̽�|a]�4�4sI6 ��t���ߨޑH:iV�0�p̛��F�����c�+�>(��zO](֧N��B 52d"N��&���CTW��&����b9݇�5Y\�%|%�|�*����ݶ����]V�)b���� Y��Țx�j��U��:�r����ـn R)Q���$^d��̔<���P{�Zf.*���G��Ӭ��1��������z���
tC�6�O|�
W�f3��c�D�����\�d���@:�۰1��ⷩb4���h�
��0q�V;
���uNkOV�m���dq���-��k�<75��<-�H��V����J�lUEMRx�)�~o��+m������s�����,��HȆ�s�}�!��w�����;b6��Y1����r��ѧu�aEO�g3�֦��[v6�p�X�x��uǩS��F�a��T��ȷ����3�E:"��2W��S���*Û���>�x���$�"5�T���'�'�i��y���%]��ga�>�G<4����<�9�@43���	��J�:���<�o�yH������Q���<��'^[�J�W�n���VѐE�Q��_oIҸH=�@��V�=>���}qI"8�n�)��6��{��y�g>�����/g@���58�#�K�p�� L�$�
<��ǵ<��u�V���C��	���$�i�f?���V|���P����qw��I�?/�pp^��/PS{�C�p ~�xpab
7E&���2z�z��s��R'j��|b������d��X�/I/x�~.�!�R�1�m��� L�л��O�l�A����x3�g���ж0�^Q#q,e������T5ص��f����>�ny��.,�>�]ƽ��z����,,��O�y\���H'�x��; ���Q���#<�%L�ƃ>��4k~kz[צ�:����P����GR�qA�����~�����5��u�n�?��vvFS8lb���_k���y�]��k� t��3�v�Ӄ9��~�������
i����]j�3�AL���S������KRʻ1�-��C��h)���z���m���2�a\����囀��y���"禬���W;�.��2\�zbV?�G߆8U)j��Z��nNJ(O�����ƌ��{\���
t�v9R�_]d���T�Hh�M]��5��Q�����{�Yz}�V>��粬17��-�*���j�Y>��J<�៮O��"�R;��DB��lI~?�/n�����'�T�Ia
��^�]Ga��vV�����%�M�ܑQ�ߔ�9���=h9�x����t����Le����C����2��i��N���{��t��a�i�V͓!����]Kʧ�(Vn��0�r	���>��f����f��'�5�g�#���|$70� a)*kl�r4�X@ז:�&�r�R�H�Tt�e��9��I�s�];Y���QK|v�C?SD�9Ե
H!���<�pJ�aʔųb*����Q���6���,4��U<���
Ά�ӯ�qҧ����s�cFE���Y:���-��������;*啧�'�c��*�"p�h]l�R@|�&��}���r���z�8��w�)�����`���M��W���מ��:$�x�π��,��rp��XO�s��&`�L�n|�(*��fU���WΠS?�a]��8���O�$���2��[���aq��-�I�# �����gE�ČS�Һ<�l)��^2G^&��y�-l���ز�-�3�]�h�
����� 	�u-��o�}�M�ѠI<���f��V�u���3��b'1~��;�����2H�/����h'��	>�p�O��V&�Im��BPZ<r�8�s��G���Y����aW+OM��={_�!PyΛ�+��^�!�lƽ�q?��	��q,co!8î�Rt���pȲ�^<6����'�y,v�1S9bh��0i+͑Ƹ�i��17��^�^����8 �:�%(C��GvqKCZ(����<iY ��S'mF��Hn�v�L�\8-��I
�t��Uto?�R\�q�	<0�����s��-J@�Jț��0��0e�Sf��^I�l�e3��Ow�L�uq��s�ڈ���xh~U ��Hvf��k�gx�Jkf����$�9�5W�ۭ�fT�J	�����O=U�xl��/����+_�y����_�u�F"��1~@G�6Ȥ7˅��'�^9O����Зf5ݾP~�m``�ƹ懵+��6l�����H����ȃ���~�|_�P�O��δ\<F<[�Ρo�5����"B^ۚj���_u�o}q���� �<<�� I�}1���i����\	p"6��L�$�=�����_(�BP
3��T����u)��>[Ai� n~��g~��F ����}���L.�^�N���`��:]F�`��2\��1v�2M���~�F3��e�j��K	a�$@�l��xt4�n^��YQ�u���8�#����r�IO��P�֝�sG*٬�^/q�Ea��������Wz��jS&��L��PB���1��n�����B����ǎ]��T��2r"�55D :s�%rB����: �'�m9�Qp�)���m�a�s�Rk@A���5���##�kF��ev��w��<7'�_=��e����̵��JR���4�h�)7U���
_w�j����%�gi`a1v�5]�+��a~lZ�.���1�.vn ֫`�b���A���<�����-]�G!�n;iKA��-T���
O�����\�7w��k�d�u���l
A��C����3Ē�q��<��m�X��2�\PCb��wa��Ea�k�˟�d{7R^p��UMs�Ō�uC'$L1�"�~m6���~�0n�s' %�6�I�y��R�~�f^x�Q�N��[�dp�.�@��ð='*�y.31�#��U����$B,�ܬ���nHa}�b���+;E�'��y�k��U��۰;Xz��J���;��lVTBbU�v�0�)���E�`48�^{��/��	f@����X��K+@����������3*�<�!�u��Cq�!��f�\d�>Yv����:�1 �6H�F(��>C߸��xÒݔ5|8l�?-朵�	�2[mF�����g�U��R\T�,���$��P�k�.���z#ƄJj���K��e?ae���޵7�����뗘?�YJ��r�:������A��g�� q�U3���Q&Za@u��{J+K�W3���[w[�[v�1��xД!��?�ƥ	���AW�R ��4�M��<�&Fh���)��~a�7�>�@r�e� 3����@j����<[$�h�;�p;g�L3�W�ns�v�/=~Q�L?�fbz��f,�L �����G�T%: BhE[�	tM�=��`,�'}�9{�Ô�&PG��u�gyq��	��'?�䂪�))�L�Z��ۈ�7�B�%�?zYZ���o}�U/�ޥor2��W27N�`	�H��p 6��]X�8A}��
���&�f�6m��7@of텄W#���^�I�ɪ�,ZU��3|n���D�G��|���R�\��8b���ш�X~�df����iY��V�F��c�$��1<����/�0۶; �n��I(@�i[/b��^n��l��U�	n�v��qR�HX�-D��v'����΂(�����|"7���i�~��K�=Z3�%����#�0��Kjc�۵(�������s���t;�Qb�\>=5u�&p!��Q����ۻJg���t��7	�_���ؓH73�"�����_Lf���5�����g��&�\~y�=\���@%+��Qh���ԍT����r��r�Z'�	ڇa|1�C� +6�,�9�E�x��Ɇu4�}��xP*��`-���!�F��8$
^�M���Z0U���kn	P�4����Lzx �r��\���NIh5��*Pd���7=t_�|=����C�4k�u^.ªD�^6P��dޜ����5UD��{vW���Ct0.�~io��0�q-T��	�tK�0S	�~�j��w)b�Y�������r}�\)�U�).H5��5 ���'�����<��\��]Md��l�}0�K��N�WU���EB�����`;\<{9�^�Ț|��μ��+R�!N�[~-ǪchԵ�+�ÔNO��}�y{|Oq��s���U�P�,�����Kq`�&�t��h�Lz����c\�*������ֿ�\�:�ƜɊ0&����6���?�ǿ4���2���0~��s����bݯ��b:�����$	��9�e���EX\n>��s���l���߁����c/�:ʨ���*b&s��گ��Bx�'H���>��p��[9�ANڧ�s����*|��w���V靁�m-/5h�S�_Z�������������3��Y؞��c\iO�t��%.<j�	��棐��!�N~�.B���������H
u{�0��?���D��:v�h��h�����3����+���;�*WB�m8n�ش��sW�w���,���ɰ���,*е�����������Z�t)_j�� <��;>n�������{�f�=h���^����A
r�و�&y���̄�y+3nq��YͰ���sPwjl&pf�&ƌ-`Qi9�(���V�����]rU����!0.�����Hkw���as�}�������~���
����z�~H:>�f:� 4u���A4Fk���廢�2�&p�ִC�@��&��V.����T��V=�c΁=���� Tp�Iz�s���T��B���a�U�B1oڢJD�6�E�~�{�dj��]���c<�.B�4�D2�:ܙ|C����k�D��Ӓ�Ь�j��d���5�>P�h���0[����1���1t��W4#(#�7ѳ�I���j��H����5ȅ3ڧ�r��4l'�o�sTh{e+z?>�I;���mt����@8ڸ�|=�w��n$ZtY���C=9T9T�e���;?�[<xp>�����6������>�Ǯc�Ǽ���X�IԮD��S�$\à2��y�����Lt'BX�/V��[��yi>�4-��$�a���еt�0�+h���ea�iY�v�͘��2��e��ݗK�����nu���MV��P��z�^S�P��e���U�^���d$����E�2�0��n\
�����c%�}ڪ?Bd�j>��-��u*�|�z�F���x寮t�m�n�<z����ܔ�k��abY�/y��u�'���\p�=��t�LI
v��A|�����|߈tēe�,".Q�\�����mj9R��MК33�8=e��ۋ��u �u@�69��v�ֺў�Ml2�?U�I��X[۞�]���~��\޻8�o�+j%9������SX��Y#}+5�1�r��鿡pz�i�o�K�;�å������4X�<S�q ��$x0��O�N�m�,ک�s� ���n�E���]��.�k���S4u�x-�|,���QW���j��z�q��m����/�nY:9)��B��O>��E�tH���G���5�^����v�3�$����е0�`��mPK�J�M���0H��k͝e( �P�F RrW%j�叝g�^˒\T�J�oU��|�zk x���{�b�
e$�G�l���?�Х&5�b���^o1�T���6o�	r��*%�ѩ�"^s#����?��>�lH�J�
-ϥ=��4�VA�MZ�}�_%II,glw c(2�3[AɎkE{�ϵ��!X����ꍚ��4�I)c�e��8�f�/�����:gD:��[$ ������q|�j$�����~�S!��g�z&X��%Ɋ0y�����'5]����������rO+P���m�Xz�b]����O�rV��Cj(�%��~R}��SU��<�8����y�����}Br����㼬|c�^������σ�l��nF��}ґ��Lk�Jt���v��T,�R�]���ע-��,��.Q~r\��N�zE��.p7bOS�d�Nab���op��
�g�R��.u��N@{.w�V�K��|��G���3Io1�F�K�f���� 2�w����uճ;,wg[�(!E����:4oN��%��� L{S�*Z/�~�U\vV�z�TRq�W�@n��|�X��9k^[;������T���t��v5����8xu�g�|���������(��39���h�kmGKz�G#�g�K���6�5��Q�_�e`/���Tڝ�{�K��E�U։�j,k�O꥓n�R�ݕ�n��M���b/��w�����y�Lt�f�0�v�&D��)k�s��Y9�����e�Y�{5M�~)Ek:�Z��Hۼk��EGELK�4_b�*n���vʗ��?�>�>��k���Z��p��j��� 3�3�n��EIP�o�]�����rf�&��k?|Շ~KT��w���-(�wŐw � �s ͖w7j x��>�ױ�A4�{�-8����F��;�_��m�P���� �{S���bV�;9�D���@�i,B$���������@=���/�1��Z�+sT�#�V�=��9&��P�K��!d��`���`͉/�X&�N:t�sa��*$�}[���L�Y<|Itj�g�k:R�z�>��bش^��>�{LM��b𦞆,���y�]	p���#�\������V�`�]h�3��)�J�^m��Y����%|�lQ`~ph�E���s������,`�ZrM�o�؉�7��?1P�%o�O%�~�B��qLy�9�@{��4z�#R��o�n;��������odC}o�Y`}�u�e��E�p��Mwu%BZ>�7F��"��A�	�I�g��(k'���؉�b}���#`}φ���|CV�����X����GX%9r 	��m}cyae�^��D	�~)�(�j.I���0M�z�����s���t�����+z�����`k�13x8��7(1=z� C� ������\��-\��n�L�3!�D���Oh��!E��FF+�Z8���s$�|���-�ǳ��+��_�\�szXª:p�ލ(ӜDn�L^U��h'6�=ظ3�7��s��[�cR��1�'T��-�k�}�us^D?l����̃Ȟ��y=�^rA��\X���G�����d�C�_�J��q5��2�h@{���=S3�k�į��ude"��-F�c<��N����}=��ET�L'Z)������S-�?
rS��eu���q�HmHm0�b=V/�D$i�"V%^��Rf'���x��7&|�P)���zt��kJ�������BO������k2�N�=b�M�>ڊ�^�>���N.����)��?�v�X�����}x<\�Z�ų�م5��("|��<��]�W�\_��>�?կE���>��K^�p�~��s\�����'쿩�N����f��o��?�s��+A���7��˛\�y<�Fm�D�����C� %Z�n�M�oN<�/���S�w��V�f�Y*����+�J��R�i}\��5vy�w5v��.��+�*I�]NSz��<�=�o>� �3� �N�{y��o1v���?qA<D�{��oz��O(ټ�^��x��Gv��]�Ҳ"6���zQ�����8kZKng׿h��� s�"]�"�Nƕ���@d?��s�XN4k�f�L��dS0��MĮ?�âƮ�3���)���wޓ�M��k��S&ث�b+z�O2TgVڑ�k���E��/��̓>���iܱo ��h����C����Q���4_w���g�&����哱��]�M��<n�w',&U+�R��<��L'/e,���r��0���W����ȑ"��(淮>��|\���=�
�*���38j�sB-���S��t��ﻒ�q� �ry<�ں���O��Y�-�����_v� ?>q����ɿ�=Bd�}�����x=��˻�HV��LI�˵���[J�*ꯎ�Ν�%��/@j�ݪ�C��욣n��V/'���VO�kݤ��9	z�b�%�>�U�~����|���Zn���!AW��P����XPK�Vޏ�֝���o�',Pԍfb!l����Md���`m�U�q��~�3��2����ГyQg%dI��K�bD��c������K�co�]kK�t���6�%��c�uiA���M/ [�O�? w���k�j�v��N����!X��?��;)�C��I�;����P�m��st�rPBŌ�Y-�j����Da{�u�Pl��"��e�Sx�9��Ҷ��qN�<�l�S���������� ��ui���Y#jξ$����<��=<�s;ŉ$wF|f��
��vy�^I��کRg���+�Q���,g{���Ȟ@�¢>���p\r�\�P<���D����(��U�x�~��pB9v�e=�_�E��=N+oNd3���~�n5qX��=Q�dX�ߺ�0q�^\2�xe�f3˼�����k����c�_�E���k��x!�g�S��Muf���W�{��:'@I������M���3�JE���h�� e3o�:-��e�֣�<��]Mo�7���;�X0�ҝ��{1��0�6(u�;f��w�l��I(��^�/X/�Ž�.�%6 �������}D�.�*�f��5��h�R��I��yM��g*�����n�m��#�oD2IT�U��sI��n�~�]g�|Q7e%�!�ecď�)���Z�v�����bA�Zo�QW�$-[\��Ri"\?�;�Gֈ��z,Ɋ��͊J>Ⱦ�_�^P�~���)������o.�=�=��b��=��1yK6?�xw���|P�P+t��x0��L2�C|jIR���O��~L[8�(��S���WR��vJW�d���)���>��:�-c��*C�դ�~t4�ypS�}�mô�֫C�}D��f�M	,�A��i��߄��{.��;�<��M��RwI3Wg˳3��Uǧ-�_�θߞn����6�G  m��mzI��:�����T���Gc�s+�R������O�N+��3�݃ė����,�\fJ����
��/.ү;ާ�$E�y\e��0����C�V�33yWw���G݇>�<֎SO��������2쮶k�5���;�s8h�����qϧ��P$�h���K�&~ا6�o��}6�_*,����L�ox������W�s�9�|��~�Nׯ#����	�����S�CrD�9l�Vg���ƶ;��M��6Qt���}*y�>:t*`���y�������k&�1y��+�ɟ�ra%�W�Q�xw#
�V��F����2r^�|���0�ٿO�p�ޛM:uS��O�Y�|��N�>;A|=.���}O��­!
��WT�}�}�#~dXYg6�����U�I7�xf���.(�ң�N��KN��H;�O�c�����*ʵ���%�s�pܞ�^���F鹤�_���j�#�4�kd�bk�SE]��_����.��|tY�oDڂ�!�a�%����e%����@��7��!澑� m{���,�"�4���!�}S�m��k.{�a��멱o{v?��>��n9͑�t��gwM�<ӬU�ҩ��5�f�M�V�S�詗b��� p阮�)B�c�� �#��o�(��A��
t�Ah�=�H��:1�e���c���I��`�z�s�Tj��лq
�["g��Nӝ9�4�?X٤�i3��Rw����\A���3͡�A���蘟K�J�7�!t3E2��N�����Հ�j�U���_K��A�o�Z*�]�w�팷</}�4B$���ȗ�O�3_�l����r��H��[Qo����ʣ:��s�rԠ���1]�mO�ʹӾ����w���"�w�+���1[6�0{6Uѯݷ��l��F}�"�����u�Wc�9��vR�N5L޶m���|Vin7<,��j2�gq��%n�ה�\�,h��i�����W7��Vf��������T��g��M�_�Z�m���XX�jY�][�u�q;��b�����]>ЋT���i3a)��;�������N����?��H���	�_=+��\�x�s��he���=H艐������jz�SO��_,]�fv	�4�kߐZ:K��O��
�����K�ג[�З�;D+	�py�ֹ�7ޥh�{����W��k8
�8f��|���B��g �-3`I�}��+�ǚj�/��ه�e_�� �i[6���CG����d��m7'd�U��=Hcy�DjH�녓����sǩ�ͧ~ޅ�s��C�G.4��\mtE��<��N�!�ͨ���e�B*}���Z����j`�9����W����lھ�纣��-�@)s�t��Tȵ�1,c�q;c����ƻ���oT�#�+~y>���s<U�5��bH�4�B���̗�����zJt$�̠�ǺeEe���0.�BY�:��Q���	�+�W�5\�	��Ӛ�q%��T)�l�{�w�2
��&�2$��G:��O���IQ��]�A�'N��k�>�K��v����#'Fu��w�l�l>4�@���G���d�2��p⪏�f }3P�Ҕ^1�/\h�qK� ��JK����
�h�Gsx�����{h5�E���Ze����ƹ�(*�(��ve�	v�[���Uɡ��ՠ@[\���D���m1�]�ł��P�������*H|�Fi*؜*��l9xV5u�*�����X��q��}m��Ǔn��ꚫ5�]��{q�c�u�`�A@
˰�R��%�V����`�Mk`�������g�(3K��,��z�#�]�k�]q�jN.��  k��{.�yX~@���{�V�~���TM�k��Q�������*�O	}��e>��������5�׭�}u��Uϥ��mD�#�-��ۗ�K�sĦV>�� MS�~Z1�-Q�XqfGc�ņBN9��Ɯ�q����҇�|1wn��r�+oG<������Q��П]s�y�냱7̞w��^:M�s4��}͸��)�hv�- (�g�I�C�W�ca���4e�a��H�y���y��W]B_z�JS�Lt�0�2�iD�j�Qe�@l��9iĪ������X��X�&l�@�U�j-4G�4@���ŧ����5��#�l�ab����6�&��@���Ӹ\�A#{[��dȤ����N����X��0\-�_�Dg�f�;ʮ?�ɴo�+�3bί�����O�ʘ����;�=k�JJw�+�ܧC\?|�D%	���ì�!���R��f�gg��c�I�(z��!��a3�~������CBP:���O8��߀�����x9o�DJ!�9���҄ �v�jQ��~K���� �9C*BN����1��T��A�G`=�DXXߌ\�ܧLϸ����gV���ٳ��z��f��P����R����&��v�G&{��0��ܫ�ҳ0(��ЯqI����c�N=&,[Un�N���ŧ�un6ɸ�v~� ��.z^���5�(_1裮��[�����/�}Y�T}q����7�Z�
4U�~��wV~*� $�Va��gz����i���� 8��^�S�*��(�oFs+Zo\�n
�p����r8��&�YJ��E�U�,���4�,#B��Y�W��Ї߲"�~B��� AVw��G����<uq*}߼�K��]\����+�5��k��S����|�W͚Ф��,y˙��z���;�`�l�ѓ�=�N��f]<�G�皛�昔������P�ͫ�v����������~�������I��W]�&%��շc���J0�y�x�q�kǎS�?����ڏ�9��Y(U6}��"6�Q���^I7��d������	��uגV�Շ��dS����?f�j	�|w]�5�*�u���N~��q��q��jEOJ��,��O�L���SSm@df��������΅�t��_��3��RR�x}{C�+��'p��z�hI�+E|����f���m��śm�
i`] +L.�-�Y�
Km����y��F�g�l�qmEI8G����ʽ�u8��aؔÌ�NY�\��Wrι}i;��]�zJ��V���e��|d-�0��Ӌͭ:H��1 ��Y_����r��}+A�4�5Ǔ꣄�D�o#TkC����a���97�� �k�S�g6�<��<E��#+zs*�h�c��K��qz��l�jz�?o���R��<O,A�ʿ|z���B��ԟ[6ƵG����7�^����^x�y��~���OL��u� �ص�ʗ����[�f���n?=AE{���i�
ǩF�3x�@���H��92h�;�7r���� ڀ����_1La�U���\���<��g3���ʊ�����.�_��;e�Ǯ&�S=�P�	;@x�����&m�lO���5[)#��i@q,�u�s�rUVf��,�hS=���	%�X�B_��s��g\�}�k	?@e)T�P�����MRi�T�J�	Tm��_�*�HAs?`����?��t�C_-��:G\,�O��x/���}�$�TmDdO�$[Z�d���e��/m����6do�1�Id��
)3�$�=C�y����������}��r.�y�uA����B5
� y)}����i���w܃�Y���\�G��L���)aW?~L>C�� �.�R2�3�I�A��/�?����J�e�pϳ"'C��
#;̾G���6Tb/$�7y(���11" y�8B��r��ur��5��&X�����7&�����"~�x��?�%�m����I��e����U���C"h^�Һ|F0D��pa��J��ś<�F�͜[T,X|�V���ִ��Jb긟z��E �\}��Sǧ��@��)Z]�.��ҷ�g�?����5� )0^t
�E���a�vs�1}頓
#b��#�&��'*v�1�C�$98�o�"�,��(j����Ew���\#��/GIɏ�x"�x	��J7D�X�A¾�	����7��X،�i@�<�t���
�Uf�!�T:�~�r�<��l_i�J���Y�y���񽮡�����K2�	� W�58)w�2K?�TrCGT;F��_kg���'������{_������9&�?`��2-�����ѣ��>#%K�5�̓�*U��DU�s�A�߅HĽ�i�-���`�̿�%�?����7'�53�}�lؘW�ܮR�	�����s0c���W~�'�}�����؎�Y#5w���=n%L���fD>�ួf��x|��?Q����&Qs(e'��q��)��g�?Ǚ����W�w��{��0�q$2������u��:X�b�Z���L��O�t���-d��/Ί���J2��P_��x-��o�(��\6��L�S�h;nR�,^X|D|�����=J~'.�7l�������;��1�]�>���$;dum1,_BQ����&.�Ç��99�N̅�p^_������i�VRH���}���r��y��M�Y۔Ͼ~n�/)����s�|��ᘾa��Ř����5�������6��oM��������D>0�ܢh�2��*,>�<���{�m\�Ќ��cYy���I�?{��i|���A����W�ʜ/)�A�dp�,�(�H����I��22�[��t��3��	-��BDSs�Y���&��p�;ϡ�8Ifz"T��=�?vο��J�9�PN�,�L?2����!3y��~(2���I���x���:y���cͰ���G�v��p���1$_m���:��Ș�cH�h�m�X~��;����N,���^���{�����E<�М�G��S��yg�Z��.=i��
��L�ID�.�T���u���������q]�fP!�.���ݪ�L�����ᎏ�X��&��RZ璎אVX��;)�c0�4�:�3ȫ�d��ԚS�����h'�rxsV�2�c������g���~S�J�J�sN�Cǧfe�����G�]��>�'��V����<QC�h�����xQ���,��i���`с���K�Y�#�ⲋ�j�rnͮ�Q��-��q���g��տ�Z��|�P�xb���̧��Wy��f;[mn1o$��%bI��(�oh����tëE�-V�E����i�{�ah��q�q��6m`�I��JGk$^�m�<��Zݖ�P����<5��߻ "�#(9%_��U�ԄN����֣4�4�c��W�Ӭ�C��/�h3o9�����vyq/^C�>1�@�@�1ʘdkP��l9�B]i8׵�`���Ϗl~jِ�H�f���G�ĆL���&j�,��������]ks�%������}�Y��R��R���$A^�Ĥ/#�w<��?J���[6q��(CMp��iL��$���n��*��i�J��s��e�jߞ\���t8��R�C�p�)�0�8;|@1@y-L�o���RMwVyl0T��S@#�_H{�W(����vj\�����@���9"?\0�E�c&#��ɀ��"c� �c�V���g�C�k*�e��k�2��롖��U���L��#��S��.Tr#-Љ����;T*G7�q���h���4B|G�'�3A[�3��
 �۩$�P�fs��P�F%�c�F�*g���*lm�{yWYD-v�Va�i�V���H��D�9M�S2���ma�AUS�6E��}��Q�Ұ��w��o��{1�6��g����8�=nHU9��X5��#�>@��2��z%�I8��M��Zb�Gz�0��$��rʂ���/��'�
<"p��A�[4�Z��:5hΦd�-���DYO����J�������*ؼ������(��Q�_������y�Sz�R���V�p׀9���k<|��4�"h�k��M/�4�(�@�&~Y����O����o����Ro-�R�oޣr>�W;������}�cZ�ػ�cK1�Bk��΀.`Q���^�|^i�D�h.�O��Q�r���&�W��K�ťñ_��"�? ���OQ�A�?��^sG[�`�4e��k4�nr@Ki���X��3��X���z��7��V�gS�Zm9%��ww�m
��$��e�4K�Hy�*���+m"~�e l0%��եg�Nr�����Ш7����`�(1�E%=
�:�ȣ/��������W7 �Bz͒J{�����y�u	C_���"�"�R�@�[�	A
�w?ү��1�L�k��8d���ҋ?��#:MY�ɘ�m�o�p�3���R��MQ�B�P�m��������/��mT<0Պ?	
&[��ra��1D�}4yA��F�;>ޜNG�L|wً�R�*C֚p��b��:��:���a��tGC��Y�u-;�~ES�r+�k��~�~u�^R���.Y�弱;�d��z�kJ����!7�m�;eA:H7�V�R6DGt�UI�~�Ak+4�t �!s�V���<߿~
BTNk\E�)B�y���`Q�Ɵ�w���.�];p���/��d�~Vq��G��w��Z���/��|�$|�H��I4l"qm=S� �[�'���h���EQ�ˀQ��=J�P��~E�#�T,ֵ5Yե/%3�p�BAm���#�׈{�y���؀�FM# �ُ���2�%˷��K��.��!��K�o˺��wo�dd�nE��{�ES�3�6�}�k��Gy-
����L��.�[\��j&@���$�V���+(%�&5)�N�?Y4���.}:�Ig�i�YW7��B�A�����H�m���_Wp�n��Su"d��M 6�" /���j���`��#�f�
}���I��c��y�L?2�d��@P���s������{�����D�����S�y��ĭ���C��Ȧ �:�
�*tx�ig戼PђPfǭ�yOP�O
[sY��:��AQ�OO��?*�w��C�B1���_z���v�m)�A�Rf_�3k�mPd���n�l����RY��/��ۈg<դ;o�~��{�u����5���#���4nfm��� ���?wɉ,
�_g����|#�қI˽q arH[Ҩw���u%;�˟�?�d)�D
�x���l��Ϥ�ӉD[$-O�<�TZ�P�S�0Ѻ�u��m�J�-sl�}�0������FL�HU���e�Κ}Z�r��k�潎 ��윭*s�o�����r@8����	���̐N��J,������F(�e�I\�l��J]��>2���^v��5�G�˼C�^�x9B��4>W_�o�'Ʈ�W|3E�pUG>�(D�f��}I����zC�y�B���ݝ��d5݊��w2v'v?�8�t�{r+]�)��Qi�����e�����$����O=���P)�=� D.X҂g^B��O(��>z���6 � �h�bI\�.��0��! Dj�y� )<���G���.�U_2�#�n�h�m�_xx
���}��Pwb�s��TB��"�ތ��O\���r[����-������l�A\���@S���Kby�3�ǔ��R��}g�Y��_$�X2��
~�{K�SX���H��Q������a,S��Z�C[��Ѡ۹�Ы��X��G��IU�[ގ�ëG��η���f��N�e=������J֣�� L��2�����WY��i!���.��頚9�l�cIfs$�C�iK��$����Dqm��Ti�JC����	XI~�����4-��hM����*�3F^���鳪j��ԍ��}Z��{��z	�	�7r/��B5A�e�T#[��9�;O��A��\�K:���IY��b��#ia�#��@=۬���
y�,�+�v'%��D`GB��j$��+A۾�b�U�!&�FϨ�@��`���o\F����G���
��#�#`bV�{̀<錡Nq��Yn�I5�k��Bh��1�[��*�'�p�;�+Iˁ�h���qܷ{FXq�!��L6�V"�h��9��T�^)m#حY@Mɻ(J����� ��`{)�M�P}3��I�Иl���`�K����Kԧe��%+v+G8_G@��,V}���{;Lav�������h����{Eam�������UEPΧ�����M��}���f�(Q��f���,u�҉I)"�X`>"\L\iT��f�jVd�uٝ��SE�'�&�,�2�_�$������Y��_ū�T�Ŭϔ**��}/�Gڷm�
���#��_��G?!=���V�Fn��k���8U�z��Ncݱw�͆�nf\�D�/7ݞ���g�����6|Œ�rz�������i�!�,"����'
�"��A�KĤPXO��pL�:і؊������v�#�щ���f��-vi;���܊f'��2����U*Pi�I��C��JGZ��I��Y��z���T9���H.�+uW:�M��'����5_ @��уG!k�n@uuY}�F��X0�##�a��%��^R{��c��د����O�i�-�:c�t�tE��j'��ZT��v+��f�BN5�����G"����Ybl
h+4I9�O��K9�
/�j��Dv��~7�	�~~i�-�}�q=�)M���q��Sv�Ԃ�����)�0�͗d6E�=���2	�jV�r�G�C��Jh<��J
A�\O����d+�C�H����r����=�ۀA;b:EL�k����wW����<VyF�d]�,��T�N��$3� j�b���c饊��W�",u'L�,���!�V���%��[�h
��U��hA[j�|Om�K��.�������ߑ��eA�wf�J�v�k9�x��>�g� _X����d���I��x�h�}�.hKy5�}0�?�����"`�	9H[���L�e�c�ƚ���	�7�ZG##\}�\�E��(B����_���ؚ�ZX� ���ׂ{c��&
kQ���:Ơ����hSC��	�Ǐ��@��"�����#�m�_�1`��oAz��·���z�~F�̗�N��\9u��Ga�Cm;�o;Ѳ���J"pʯ.�R���co�!���]\۩��<���+�o�}P+KB'V<�QP7f�a-iE0Č/P~�r��:�EHQ��gУjش�<�w�#�~��>�2�#ϺϦӏ⪡�����8�<���IZ���� �KC���n~�CJ����(�{�zr��6k�F��<S�8ѫ����������_�o%H����� $�a������=n��||Y�rӹ6s>�9r�����h�ͦ1NaUc�^����T��)�g������ (�T�F1_�,�+���"�6�Tٮ>�z�r	h�d`�Fe���Z�������� k=& �l*._�͡��V�qy�����pv��nE)?�����\�*��ꎽ]SI�y=�6�7$��5iq����CO��$.z�UJ���.X���u��7>߰��m�kW�J�"D1����ؽ��nV�x �5g������l&����+1�s������[9���I݀\z���:�ɮ����o4D[2��%�"\���V�>$"V��nFh�)���+�9@`k�5�Q���[���8��L�7w�v�F��9����!���?���I2�����9>�_)3��Q.g7�������5U����˝ή��ƼM8�>�A�7�]�[ȭ�C���dy� �t�lP�����x#�,���l�A!IpXˌf}>[WgL�q�0�7Ra|q����6��nL�K9�$N��sY�;�Kc �C�!� z�B�E|��kH���h��;?�%���8�L��;�T��a!ҳ�-6��>�|Cŵ���z.:�z�T0d�j�ǯ�?�!�����J:�J�𮕨B}��0E	.��Z�ibLA�=��X��X����FR����Ur�K�90n:���S����:�f���%_��)���+D�|G�p��RZ��'�*��3W3�h9�R	��/؈���!��]�l���TÐ.�>�h�	����4B��Y��4���+�B����br����ElH�xM�N�f��9!��TU���9F&�*�o�m�΄�ܐv4�Hs�����?<\���6G~W�����}wN�nv��h퉇b^���S����U�}�$q�X=��ʙ&C�=���#&h��^�J��J�ω{j��2,��k���Ŕi	�]�p=4�[�t���sf��!<���2���=��1e/�B�+�m�iYm#�j��;ڢM�M �Mh=��˺����Ha3U�)b�OϞ�+,<��Y��̓w9_�*DRU�翨�1@�D��O/�k��e��s����޺e,�!-��4�ިN�����]�G�pM�$���(b�}�Gv��vy�����S�U˃ՙ��> �_����6��k��vc3�1�:��ɫW��Z��VP�hJ-��6����J���/�@	��C-T�"-3A��W�@��E=RE�fFQ3a��.���t"p���j�P�8�O���F��:F�J�RM	y����b��=Q�d!��·��}��L�>�o�ӧ4b�*��zUd-W���S�&���ཡ��}� �ĵߧ�/zE;�F�5�r�%u������G���ɸ�窣y�Y�u��o����Û1�7r!��y��N������v�X�'8�����P��L��Íd1��A���Sc"ugk}G;�[	,%�����e\)�~#���E���ɠy|=�^�k/7�#���kP�n�J��/�b�sP����"�NSS
��H�Bٻ�aF���4�f#�g��]���������	�=�&v�!����Oߙv���܋�أ�}b٣u�;7=p��8�RF雷{����
-���	����=ֵ)#��7�YH������ L�n3�I�z��$!A}���](��k������D	����^�1Nj�Ԕ��_X�.��9�����&f������E����(5ID
�l��N����܌���YX�8��	(�a�~�8Ŧ�D�+/��{?���	T����D�G��7S�
�S�g�*+�2�EX�L7Vl��1�&�N��qc6Ux��X�#
Gc^i⯢�̠�iv`�}"F��!s�%��q�Kby��+��~���"iL�Z���j�/&�3��s_̉�����+'���'���/�ld��ȡ ��c�����cjJ0L#��>����O-p�6�>���T�-�\��P��y��n���x�Wc{�1t�q���Vl��nw�. v�D\�cG>a��I�`�鵋.�������@��A�P����>�%s{�E�܄�����;u�/�"nA���W0|,%c:ח[ƺL�tD�p6����^ ��0Wo�� �U{-n����`gv����}���Ӓ��jr	��s�}Ox�&�vc�	�#�#`Wq����ݍ�-�����h�"'��^��I���{8�d�r5hz��M�H�s!�cP�l틉w����y�Mc�����v�+GA����8�n��!?v>�,i��f�#'˜@���{�[�j���3�8�Q�.��Zn0�|E�Q����ƾ����U��-Tax ��	��K�O�O5�^�7��L�o��m�����1���y��s��<�$�33�UKG����4��q#iU��d�Y�G�N���5�7��v�ܧ
s��S"l[�� [!}n�$��`�P��@��9�u�{��[(����DP�h����)��TW��o����崒h�3;��Q�o��pK� [~0�a���eW�d�c� ��<l
ɮ�H �߽�vH����ʎ��@l�v�49T��S�.2�P�u�{J�d��E��k�c�&9G�,)����DUzW W�o����P<Õ��x��%XL�K矃[`���lvbw\a�'�Bo�z�;��qh>F�%>�U��\.�(�jA�߃X���d�`���O�Ebp�5b���'�!�-v�un��V4��՚1�����Bkqb�D���P���
�Vj��Kw"2�	`3��g�Hb9�+GL:c�Y����W�M$B��"��%�.r"�J��V#|m�a��Ƒ/�u:�Zas ����Ɨ�x���?����WIY2�(-g���Ҹ&�w�-4�]����p�>���a���Ԝ g!'�	�yZ?��P;xMea3�)�ȶ����,�����l�N,<w������� ��ȥ\}+���o���0H�3uP|]��pA>�������1�M��kG��y�v�)b/u^v+BX����sS}�������� �zz"R�ZnU�P|��]�b��J��&d��#��>�ɣ]��1%�y8��e�_%;H}i��>l�K�.���.�|{ ��]8d,�Ѡ��-#	���.�{���U�A#���=�R3 ��5�
C�q�zJ�ѭahr|���MD�=�9�M����FA�ĝ+�c��n��ޕ�����b�v.ԧx�*���S�u��\5=�<�ZCY��j�y�t��y!!�X]��,�f�[�������wy����u��?����H�g�q�S&���:�� � g�|��0��G�#��U�V��OQ|��L��o�FڏD�v��S���;�3c�~N3C�ȥA�cf�P�	����P�t�� ���q�g%�\��ZW{�3I	�ȸ�������4�P�!���[@�U@���$��|��w�Xz/x�6r�����C3i�\�U��	�Ud�([� �6 ��B�w�m�Vt�pP���K�� �V L������B�B�K��Ԫ)AׇU�O��>����'����FҾ��g'x��j���
i�{(��Bw�[�'8��MQHp�UX�`!��g��)�	��9�Q:1;�<f�8r�c\ ���CN�||ǜbW�$0!R��?I����v���K^�ٗm����}ƾb�-'�z�ȑ��8�Ya ��_oj
ő�l>��b���Y|WU�3���R0�E]X�ϟ�"��������B����s�ϓt�]Q�� 6�'WTj�D��3��l�щ��k�����������#ha�����Į
��mWb���9�Q}��K�~����Gȃډ"U��	�:H�Bu7���z� {�8천�*�}|u��Ò�ͨ��7eVF8�<�"�Ŧ�Դ�2��aL�lщ R��g�|qD�۬����(Q����S}|�����3���]F�?!=�o *'3��B���?�C?���JU��Fƾ"��J��l�%���<ZL!^�����M?&���}��� ����9��m�g�n�3�7&c3-'K����#�����)� �O���oY�s�؍�)cɾ��*�W!x9�y�����͘s�j�ܟ9��Fe[ִ�ϧ��&��c=���3GVJ���5���_�7�п�'�\���:�LLM-�<<|��g����lWP[N$o��
�"ѥV���4,^:A�Id�j�d�U�	�EQ�u��=�(� ]p�l���2��
�w���58���>�H���-���Ү�q��6�K�`�Z��GY�;��oh�O͢}��.�P/˔��|0P�ڒ�)��}�;�%�L�N!ץ��&\rz��W=�㓞�i��m����Y5���5>r�MF�p�l��vR�v��_V�Y.�\�盈���
f\Y��X
A-�j�O�u+�#���c�5,�C}�������Wz>O�0���ֶ:��I�O;��j�a9�.+2���{\�n9i_��������č�:�y��荙Qsu�>-��1˥ɥ�Tn�J �q���VTm�����Y7��jB���}���+`��z-�+���R4r�&�F׌(y�H���{Y�&ǩ�# ���U$9%��#O��z���鲠WlQ;���CQ����ݒ��3�V��������r�{��p��w����$���5�!Vw͋�r�Fk[7���/�P�GɽK)�pn�Uk�(��<^�0x�J�7\B^2����.��Y��WA^�}Ц2>�����ݛ<�v��@6a��5F,�%�SE��b������h�j[,6�o��K䝵s��˃��?��/��� ����� �&�=�RSDG��%k��-��\wY���;d�P���`Ä�B$W��U(?���P�0P̈���Ѽ޿4��ޏ<|S���QMs�Zz
jO����	E�g3�I�G+#Uk����*��o\�.�m�T�u��u��27h��~4��8��8�-Z��8�#�'���=��q�W���y�m�z��a�K�_���Kmg,�m;T�e��f
f;�m��z`�ti��j�TC�O��E�C�?�c�Z�LP�o�$X3 ir$���_�BG�����&��Y���S������m�a�HC�M��<~X�w��^�#��[~����q�j�ɪX�{��1���h���O�N�+����q�ht�3@G�SYC*��-��vz�����nٚޱ�O��	��Jx{A��,gk���#}����9f���׋s���X�(��A�pZ�X����PK   6��XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   6��XF���?� Q� /   images/f590943e-678c-44eb-a174-3243ba5f3820.pngl|	<Tk���ܴ*�})�F)�2�t�d�2�L������'�m�si,Y��kBc�Pѐe�C��4&��4���ֽ��}���u�s��[����9�~�і��!��sdS%"�^��I�J�<��}���z�߽�7���7x��BC ����V5:_6(�ex����������__�C�n(��u�C�w�Rg�d!��c�?/��}Ƥ�X�P�#�}�`bVO-NX>��)��l��T�z?Jo���c�!P����[zl����e�Kyĥ��j�������v(~9�9�D�FWo5�`�~NA�L�L�4�M���-;:�6RT��!f�Y� "��!ɱ�����?�snRr�D��n:��8���0Y�T�Ip��Ҝ�Q�A�-f.u<��}��Ha9�:�C#J?~��X��s&�D�W��t|�ljt�X�g���x<�K_�C�LV�},�2�����Yw�揹ճ�<	WF�x��C4[K�9�p��8�愝���c������4r�3�v�R����X����i`O���-��LȊ���G��	H������hhiu�r�ׯ_37lےlY���~�Z4d�6�I�革��)%�ͩ�Q�[MF�)�OV��n0��X3<S�/}K�M�8hD�2Ϟ��s������ ����~G
+���i�j�[ZZ�c�cta���{ZJ֡.�����m��cɵG?�Zpm���k�����9ׯ>q��U�X�Y�P���Y����_P5��a*���z�$LT偽��;4Hè�<H�(�?�t2��s��;f�9w�O!U7��b�+]�){1K� ��"[]�c�d�z�0Oa�[����s�>���2(�|�z��[�?�����
K�9n���&�J�����Q:���rrrF�
�^�0y���ݾ��P�8�is/3���CE\b�m�7��'���%젡A�֝��)n�;o$�)Y�?cd4�����ǲ�W���4�+���H�V8J�&55�iek��	-iӥ��PW��*��CCz~�G_7Źn�s�_w��G�m��ϋ~�U�dkih�KjC�]1� ̈W��0�펻�Mx��������$M���-L���{�����u�B>�~�Z��"T�>11�+�������В��8���B����l�C�:4���y�;�W�$#<�$�����S�z~�"2i>5v���Є����� =���h�[߄ɓQ(��	�o}��*Q�=�9�"�V���� �*�6�^�V��k����:LY�Pc31�qP,�«�gZ�����V�vЈ��$�1؂�|�]4z�`'�mB�w�F=��[vo��0�����\�����@������m�W����ю�g|S���q��f?��p��5 3C�_��+�'�R�?���Y�S����GLE�����	Ӡw��qa�d..�\�z;�m�:==m�����4)g*�*1�d�a��������'�-F\�	[����;����k����!�,l|t��b^�z�����*��+[w�ҕ��Slg����	c���or����Z�$�*
��@�����mq��jPG��5 ������K��}��v��q�X�=a7Ƀ���g���C�>k�Mi[������z���$���wk�Υ䌔�|�����Q��w���9S�z
79�8W��7�<����ٗ�fh7kM���0��X�>���3҂�<�B)��֋ZK��uF>&�<�2-hjjZ�|��T����-�2���!�xF���K4즕O8:&|Yp���S�{j�2���t�J�0�'���5�ZwX>��_�/P��3;t7��co�ȉ�Ŝ1��C#T��I��N-����k(�KR�
�:y�q��9�N!�.?���s� ��j��L�b9��&����?b���*d�C4�ew�nU`$aAE�x�n��2e�J4%!�d�.������8	�MCVBP�!���f�U��#�g)�s�]: ��������chu�u�(#X�R�h��M	�%�Ȭ��HE���J�٤<�,�#��B(Uc�̗mo�r!(��	�'�s��I���`��BBQ�K�[GS�dՍ�
(�C�ְ�n��m�n;4�JZ���|٢��i�]V"�':��-�����|K�s@��'��` ٿ�A�k
��~��^
+[RJ*���c� ks�vxpQL�� ����&��4"��Lb�%���	��w�`��i�r��
��"S����-hw�5
��B� �x��՘�b薞��;�(_8�\z��z7 �\����u];#�U#�ΊYY���Oꅄ]�������N�n�.]�!k�ϤZY3�@X��ϰ*9�	���Z9%wd-��m�C[;�Vi	��gR9��YX��1AŘr2�k����I�e�oL�c�c X�� �$��I�-Q��3��`8	YP�UsA��O/o�)hn��]����H��y�H*沠���G�F�'�b�U�<HýN��z�{y�ʕ�/kk���.U�iC��N�e���lmm�}H:L�W�jF����I��u|�OB�*�%g	\N�m��vL�e�Ӷ��I�A�4�����_L/C�I�h�9F���*56�!�UyO,Uc�P�r&MQ�e��5��s�TM�AAW����w�+=�ב�5�I�>UNva���v���������%:2ק;t�$1yX��w'�7��9dڥ������,��ij���dV��?�*Q�B���`�3~#�	�/�#I5AE=.#�}�W!f'a�9���Y����~w�"(_K���Q��
�
햘��2{ s�M-x�.X���%R�NN`Q��,�Ȭ���%�K�U�xʣ{����o�?|�y���Y���Xe��ή���a�3�P�|:)_�T�8:�<�����%VUa�����ci�������ɒ^��ީHP.��=��WJ�����,w�()��
HWu�c�&d�=Z�ܢ��V���~�
g�HR�����J�u(���5����#Y�*��V����g�����h-�4�͛7�C�x��m��w
����^����~��Et�̉�A�P𷾒�T��״��)~ޚ~�7ԃף�W΂��HU�����\`�ϸ�Z�s:��Y4]p��H���q�o			�Qw���q�� د�`u���O~d��2���hJ}�x_x��V*��xcE�O� m-����f��1��\z�[�a���5~���q��
�~���7W��i͚#?���t[�74|q�ҴO�~--U��~�t@Q�5�5J�^�Ч�%���A�Z\Π2�[l0Ӫ���d�_��ͥ[T?/{�CXy��d:>U�-	l�"[)w�#�Ȕ�4\&�Zv��GJ��>ё�Z94�7�ݯhJ3���$O���m꟡�K�$�Q_��Rą&$�R�U;�$vu*���Sæ�g\,������,G�.����ڵ1�S��T-��K��j�#\�����]-�E?�E��a8��C��N�[1�ND&k��M�R-���ʺ^1� R�\)������oʂF  �W�1Z�����Q쨿i�P N3�S8%a*��L�f_r~V�b�+��^��G�PO[ͬ�W�k^�0��:{�R�^�?�iW��,���&�ciG0h���2N%|K���h4���{>4�Җt��C  �L�u�uu{<p�@1H\�U���_7�V�������A���w #��z�Rw��T�KR,έ3s|f�!I�_ܓO	��֥D�$YY3������41�}��OCכV���I"�a8# �G@���,�~]�:�<Y�f��ے|H��R��a.�Ӽ������TA����MK�u"9i���	CD�W��~>e���_v:�v)4�4"�'%x���CG<[E��������圲�m�»K�=���#�$ǥ`n�?�P�O��K��m���Zch��m�̅}�����U1O�"����8���.�X��/s�>����&���50R���V�ڏI�pR�&�Ӯ�y�Zk|��#U��I!�^x�f�pEo��"�!��P��@�f"ml�&�v�릓"�%��"����JZfv+�AO� ���2�a5^-W�K�C	bѝ'���.����Z�r��/ՏرI�u��&��/Țī�d��s��< x�B~�����I=j��dA#0$����Ǥ���P�)�X3���Q�����i�z��?(�u�9M΀ѩ�@M���j�#!��-��G&�dD��5S!U��s��C�$t̘�i�Q��w�_�����1W2 ��\�V@�3�f鹱R����)A���;���p�L~d��(?��%�Չ����G�6���-���p���sI � IKծ��)�U�a�j�T�{�ek� ��Y�_;t�M�Z�L���i���e3	)]A/�;|��?�P��ى��{2�H����h�n�D�00QK�Lm&w�=��� 2�~N�Z������yMj� ���٢��AX��3�OcY��G��~�F�k6=��k��-E�U1��1�맽�ۀ�ݿ��OSu�A��P����U����IU����s9@y�[X`���۩�`�Iy�x�.���=.�\gu�,u�oo7�7��=H���Q9)��p�jh�XR������)	�(�j��DS�i��:� ���j�㳚��Z�Qů�+���n}{�8顰h�}o�����5�Q��3N�GL.'~=O��*�����@%iFFizfP�>�~ke조�g)�w�7������������r���C�?,��<�:~2f\ic��+fچD��#����m��H69ZQ�Hf���}��5��G���OH#G��g���%�H�U]��SIQn��C&�pg ��D��Y��{-�~�a-��䍞�'!3@N��4 '��%���_�jN�j���D�e�_���Am�z{��LBաm<A�l>��~���w��"*=�v������QU�$2�(��cƟ�u���wg�bT��ӧ�����1�9������ 0I>�����ם���������6������3��ez��G[,����ݛ�x����q�׾(�U�[�ܡg��?M),�*�7���L�q>�c|��N���j��@ ������㒒�'%?�H|VX\�:=�2)���Jm��>��=c�w���G�4Z%�w��'�(���F��6X��M�θE=��3�M�E�ȯ�=���j��e�V�1jpn����8^��a"�Ls`7M��Z�#y��?;�~ÚS��`���*�� ._+�R��PL#�yY���JJ�~�c�����csW}�6:�� �]�*���B�Aw�E?}�o�� �Z_\W��q$�w�B�˹��n�F�Q���a
]�����։�F����WQv�9�HU�������/UT�u�LN��C�9W��%��\5_��TSY��>�/�� `^��5�wSԞ-�_�W�%Ri�vĴK���7��P�=������4�J��zr��c�E�ȇ�_ذ�/,������&D|r����^U����o�t-�-�)Y���u-�w�s[�Aީ�`�㼈Gx��م\�;f�\�3��L������ٷ���?�1��ia��y禕�0��
@�pn����Yl@��&Oyvzr�ZDV�#R��f�*��1�w���j�!r�"W+q(:A���eV@Qk-�[������.�u���$�7m4���_�1݁"�P����y�a�Zdem�7I���n�³)Z��2���4_e
	�sN�m�^�.�CjjCW�nm��+�}�h5��N�j[���凢���	a���ǫ,m���K�� ��IG�y�J c�4^E�T��ӪV{_8/�H�7:�Ǡ�<��᰷�#孩\]y��4jd7f[KI^������=ԡk�g:V������s��R��{�,�D�c�����g4�n�X�k�,B��DI�[1��,h�����D�T�נZ�2%����9��*q�N띌a�
��?��j�nYP�q�h`(3SD�"`�w,,N� QX��{��1A{(��G/m��c�xUPv	MMM����}ʇ�˟J�̎�qJ�e�`w5�p�T)��~�8����[��)��I��h��
��AӮ������[bק_���į7m�d����nN��Ҏ��tƑ�4?��'(���oOÌ����$�i^�V;Zf�>?br�'o��gB�3��'� +�]����K0)+%z황*��*Uc�$�2��i��]�I��,Ѵ#����V��F�����SD`�t5�i���ԡΌ9c�#�7�幖A��QOTtƙ�5NQ�J�9si �ʀy��Th� x9����t�aGQUj�Y���/�:H��� Ĥ|W!4"�TUᥛ��z�e���?�!!�E����30{5W���Si-=n`�ۥ3F�����9QF�{���� �8�NK�>Vk�y����ㇺ0�-ӭ~�bG�$ �:dr�4'� w�m-u����G���4\wg�8����y���>k��x�3�ǃ�@�Ք��q�w�rA��T0~Vt�Qg���6G���(��O�U�����y0!�6�ݧ��e�^�^�2)o~�U��Zм5�4Z����V�����$>:��4V
(��1)� I�H�#L�`��E�Ӈ�ڀ����^�`^aVgU_�OW�*�Jޯ�D�F"��OSo�R�[�Ј�=�v��%|�|��Vh��މ�͖5���¿"o��_$��Q���o�v��!Z7�H��S�/�h�C���G���ju�s<I6;���w�|o?iv���u��T�<m^��_ ,�\�W��f����o��"0�b$g�����6�boP4^+�Zsb�W�^��_� �?�.U��W|n~]ON��?�"&�5��j���<P�����"���K
��,<j��� �(E�aFL����yj�� ��a�C�U�s��x����M���5=3nۈDv�AЖQ��|���K�9�k5��wh!i�z\lu�v:��ȕ��Y?��l,�E��rk��w�1c<�p�T%�@\�&.���J���Ʒ��!=B��^�>=	y��42H_�[���A=���������&�
�Ne�������=��M�.�at�J�+�����q�1�w ��M�� ��y(ߢ�5iJ��М,����p��.�H�	�eC#���	n���,�W����a_8#-,�?\�-�!��U^�o�(��tȄl�������6|�I:�Z�{�b~ާ�-�`���>)CA��~I@�LB��D�������g�d�;v�lK�X���l)b�Ԥ��+`h��A~��$Ŗ����ر>�H E�
��6�8hć��.���0���ݘN�d�Ii�ޥ�cV���U�F�����K�c���E���H�M�m��a�_�}3�۰0(.�C��!�m+��!��X�v����ج�}܈_?�_��$�<���(=w��漟�E�����q�n`N�.-9a��?-�/��Z� ��3����Ɇ�.����駤 �`���U�Ӊ��*Q����%�B��-|"h``�z�h��Ќ	f�x�i�\��ޭ
����ڻ�g�c3��R�L1ݖCKZ��U=.
@�ې�Z�����A��Bb��+|�C���C�KK$
G:��h7�׷x�b0����@�i�nz�v�a[��c��?(��-S �%��(�<! y�$���A�!�����),����] n�~�����?��@V��e����.$���ƨ���Q�3W8`�g����κ�)���`O�Y?T��X KF�`6^˴ ?�v���.&&��+����^��g�ysz�n��Y��E@�2A���2�^��p�>��m*�qNZ�"��k���X�����j�E��5�OYw��U���<��@�M��f�F��Jĕ�5i�f��Cp�-�N!��4Qx%h[��2��V�?@�u�܊�%Qt��_:����=���ZXD���fA\¼���ʀ{�T�T�Ϡ.ֹ�C��}�TQ��ώV専?�=�#�3z�W4��
ű2X����h\��9JkVڡ(�{�Vx�ϊB�Vx�M[�(���x�k�β���e�0��Sk�����y��Yf5���L\�q����Ќ�h����b(���T��
���}�M
��g�+��B5��h8��	�;�q���(��Ո��ۥ{$Vim��3�N7�4	���< �C�!��c����	ߎy��G�OH;Y�3皥�����vwu�� ������8�������ɾ&�ed�<<���Mݴ�@64�"%��+�p�*Q�����6v�g��z���+UcyT�P���z@0��qr������)�P�|�< ����~�a%�l�]�ݟo�:V��D(wu�DK���Q��#�G�D���ߘM�	1Ka:w6��b���٤�VӔ�^K�g�n�0��}�����f3	o R��J�	 :«W^}ά���H�N����b�/raqtŷ�T�\KG'���Kt=�s���>�(�S��h^?��G�5'����@�]�^VU-}��7�~DAf[M�kmںv�g�Ry�����s�IRn�O�a�;"Ǆ���fE��| �@��s���7�&����sQx���� �Q�&�!1������ń�����%�H��Ɩ�}� x���DFY�ҵ�K�
��%��,������ͯ�|Y���\���a~~>��G|�Լ�e`�k%����d^P�*�6!�~���A��n}� ���r���$윙D�3^�n� Y��q�~A+8��#��`9فEXD�1�Pk���p�߰0��k�V;Dn���y�]9_D��x��G[�į�_8�Y@ht�++���s��H�+��yo���k���b2e��.�H���D)9��
��g�����!x��a�-��W! �H;�N�Cn5.�^"g��v�4�A��T�R�lm,�S��ݭo&��s�;��B)+�i1��ouEM�J8�ѿ�c�# �]����p�����cW�����u�"��7%�μ?`2s)�L>�*��=�������R k��ja���� ���{XLLX:}b"����ػʄ����9����ukd6�s�Fgܩ�H����u��/.=w<������������m�H�y�<�wU�OU�>���Xw��B�d����ŽO�*�nҭJ�9[�=����d����O_�'��\O���R���|B���"���=䪄Cn�H�L:�ʈ�v��ѣ�j���B�y�o�(i��Wl���?Y욡���<G����
h�c��Z���I��֦8���@���gzC��u�q j5�Nw�����o��Vhp�O�=�
�D�0�t�hĖo��t'n5A��^�3�)ƙ�Y�[�!����F�oO�tp��@��Y���{����}�^�J��T�s�f��A�w�F>)�
��%ԩx����^�u�����-QWlzKo60x1��\�DL,���ϻ򿳃vӐ�� V�IyWgq[di�e�?�a&zyU��mbJB�)`_i����H�O��tǅ�Һ�w����2ib�X?Xj��!{��U�W�%7�<OG�p�Ϛ�e<qMo &_X^\x��5;��O>b��0����/��m��d��'6�1#'�Y�|!��	��3!�����C�f͎��@���Oޮ��D�{�{! 6+���Kx��o��oh�ZJ6���N���6��~{�L�DV2��)�b�l���tU�����9 ���e���U���.��Pl��'�*���"�'77��V�b���_����m�	��Ժ��!A�l�"���@�7��v�wU��-�?���D�|�	����uğ��f�nB3��Kz���<N��2�f=�i��p	2��B�$��)�б�k�Tp�꟝��ֈ�����s�۫�ܤ�H��,�X�����:���]�����.ܳ��
�����"Z@�9R[^� *f�!ݹYSV�����w�?yb��z�7�wr�Ԑ��>��Gn	=�q���G��o�����>ee���+�M(Ģ�	u�H�_az/�ZG�����2�0}�\�B٧<�!��-��o{���qX�*�h�#_\�q��Rz�3�n7&7���>�+�d�
���;`���W���ߒ��-Y'�|Qػ?�o��_�g�����`M������He]݊����1H<����_bQ��ɒXe�z�:1�^�dg0�V���P��<��}L^T}s��u_�3��Fd����4s:����6JO�v��[OZ1�W&Of�Y[��{���F���~M���m8� � ���f�G�[���ɣ!�aa�nn�Z��jm�1������Cۚx�:͉O�ɛ����G�wj�;���8^�B���b��6��s��f}'�3��b:�(��LU�K>���c�x��)ͻ>wvP*�O�Lh-�~�������P& ��2nFUuJ���ʽ�9�i���ʐ<��Zf6����p��^� ���Y;�h����҈A��l�r���1զ/&i�6��6�?��8Nڠ�}���˩qW�]��J�<H�间{��ɣ��N(|���>���E�ޣ~�?:��;x���o��gk�x��vŌ|��͋.�ة��h��)mFɳ蝯���B����������7^�kK��:S�֪(�2���ܪ�|9���Mi/��?����]tyE��0��2�/e�����M��[_\��{aq������I�z��/�."v�#g�|��\Z��)�+{��ߡ{f��\��q�S��+͉�x��ZS��p����Y7#�r�.���D��� C[^43��_1�ƍ0�����7��iڀ����A�<Ԑ~�r�����ϗ@�AΈF��U�ѩED�z?М0nN. w�{ﮘ��j~��d���s-�*/�H���z�ޡ��ba�_��^��G`K�T-�B����dr)�|�X%d���T��?����3��]V�m�::1팤9����P1��;V
'Q���l7.V��	E뷓0I��Nv�}�sA��ެ3ˣU�O_5N��c�m���[g��=��˷܈��p1�ysr��_��|K��桋(�� ]>{�=������{T���ZE��E�h["�P���wȴ�P�Β>�C|
���5m�=����>5��n�/����Ϊ:�q�m�ʠ��dM.5'�J;�ǧ��y��E�=��_��{��,h�����̢��<i`{R^�.ñ^���f��X\PP��ݡ�]D��Z�V���f��}���v����^56f���.o�mT|t���{m�њR.xqN����}����t(�YV4�,f�C�4���ȇWRUu/M ��| qd��o��cR���icVAL�]�O�8|B�J�6�U�ɲu���\� ����vt��{���_�}>�O�D�G��ʵ��UF���?	���ڡ��-�МwW��D!�������'�1?:�d&��hZ���l&�kw�(�@����=����"ö(�݃��J��9��n	m���G8������S�\�瞙���seu���t�p$O���;m� ��]zܑ�������v�Z��d
�ޭ���-��$�m���0ϏD!�m����	�
_KKˑ}�rO>d�>v�s��٪ sOK^5z97q8Z3�0�"Rg���m�(�x��#�z����	;��_���6�T��Y�t��c��[�&�#�O}�7_RϿ�� ����rƚGI��m]r�m�$K�8���F���N�������"��`�	���cEG��!�5g�l4����O���,D֟(��'\A�Ū��h��,��k,�J&	r�ǎ��� )�&�_��$�\�w�9��t��g���2�˷da1KV�f(�����b�)�姞�#`*���H�e(�����W�>��?�#EG���������5.g]���zR�y���{�G�vV5�7�hX/�s�(�����kH���wke='�<�-�-C�`NH��V���o��O�w�ӌ�7��Q�\.�V�1�KK�k:�!d$� ��F��E�v��[�+r��M/����r���C�{�9�v5������n���%Χ�����L�w�{�����-��l�� �H4�@e��TW.�Y˔�:n>�����t���OٗKBC�Șb���%�t��UU:CCC���Jw�]f8ѪW��η�2'��A��2�Zz^��+�Q�CHB�mY�qѵ�U�f����7#e����i��?����0����V���1��T���OF�77�q�N� #Q�������z4znPlvP���?�z�CAJ�?2�c[8��u^�w�$Eu��������$;�j�:���hek�]��A�F8)��L��&��.f0Y�O�7Lo�1�"W)��-'��+�X��n��7��W��:9��l�v�l�{7����8�ʙ��Znl_ac;������⏒����0�G����,(�	��G,��g=�w1�(�@�`_� �A��wI��������sA��P�H62
���'L>�j��1� F}�Z+��F|���4�9�\��K�3E��O�E��U6�s��yJ6v;�N�~���zl'�����?�EC�	�� T���lI����'��7����O�\:�{�;�� ��g*�Ouv#�	W�,bg+Fh��G�%j��.�~��v�	z=)�}�LN5�g�Dz���y��ӏ6��D�������/.��r&ޙp]t��p�-|JY��q�0~2���,j�m{��n2�,�CM�Q��}�H�oq�od���\�?�����5G�i�8i�+?�:ې8$�8��ԛ��I���j��]&w��0xB"�؝�]&(������{��&]_�p?�S�)K�M�KT3`$�Vf>�[3\ lB������0ޤso;��@�0��:�Lo�Ѩ���c&!�q���|jҋ�S���N}i���Ih�ܳ �T�	*Td����>�6'�Z�V��Z���+Y�/����O�ϢEA�K��"NH@6�ʍ�U��1� ��㩝w1>rM��B�11�?LE�j�Q|�8d�WU�:$��s�	����w�S1��g�3߾��_)K/j�+rv;��,#�K�r�D�Fl��=�9�\d���O8�C��������r� }�uO ߰J����5��c*�P�Ig�j�S�(:��2�����f�O��R0������|red������՘Z�>���MȖ2(�Wߴ�>�x�:Z;lja�{�^�����_���Tp5;H���V��\S���h���I~��/r���r ��y��\��m1<�z��p��!6�|XG��U7WegC o/��D��O�?y<!E~�״gn$�H�? G�������K���EE}�QI�/Z���8����:A-�m�������܃�욒P�Y�ʙ����:appǜW�@O�I3N���B�,���$q�5n���A.m�)�a�gy�U�)I>��ᣟ�CT5H�m|t�j��{ �D�� ������օO����'���I�+�|�ĦDa��j�?^H"f�"��s۱�/�[�J�:G�,lV��T����k�G��ÌH�^*�r���{h���'�^sɞ�Y����4��R���K<s�%��V����$I�O��٧���#��	��%
��؟;?[' lM��Ӧ?)��x[[3�	�Q�u#i:Nwj��]Cic(��a��$*���R��v����A*h�Z�&H�o�$��X5��
��_k�6��`b �I��q����3��؈�{Dܗ����E���=65���)Ȍ����*VY�՜�F2SS�����ݸYU�щ)�>��*��������U~;A�����x��������IV�Q	��U�~�OD�v�$��,V�3>A��KU 3k��d�9��k\�V�Ygxۀ�!����0v�
��� �q���r�OC�.@�� 	���$$)��َVkݮ��]2h��֋�<���E��0�#{4e�:���gᰟ�B��b�V���SƽtIK=���p���M��m�����o���r��a�M��	��Ah�x�Vt���U�͸��z3�,�B=��LE^}�h���^F�iq0� �}��"��0���Ji7���v�H�R���G���׌��F�/,��-3�'`�*s�U��Տ�u*>���)!e��`]��#��d�$����!�F;)}�H	`�!d�*x̠����^��	�ʲ"X����i�jR��/�x�r�����F����=������l�x�A�<uӕ���#MӮ�s�UG���� u��%/(���I��6��T�ͣ��)FF�у��c~z�X=A�>p?�����K�1vg^���N|��]�@�)Ƃ�hl w�R�{���
<���0�y��ۍ����&��n�<�����f����3\؏�����mVe?�n�#,���ī��^�pخ��,^-P���e�oW	��.*�|���T�� ؖ��t�o� 0pb�����3B�2�W!Ig�HC�����D���' ����8�7g�}f]��n�%]��{�"�@�q��� ��7��u�8�Zj������FJ�'ϢY1��*C�n�����nK��Huτ���;y��=�MOѡb����h������}]PR.x����&�GD�\u��d��P?r�Z?��7��;y�4YY��RX���K�BpbŖ��v},=���n��$-�w�A�֧����رM�-t���i"������Ǘ����n��G�)+.�p�������{?����ɵ@W`��\Z{B�{�q1��<��������`���<� R� �V�Q?Bʨm���$���=���ksH�ݬ�����Y�(�Q@�u�Ƈj��{-�tH�Ů��`̈́�E�sJ���ᴹ����h�sJ�;���ww�`W�u�]�X<�'E�r�������0�����{�pa�4�يk�O�X��!����n�PJL
����!�9Gp?1b�[/�v�G�w�n��OF�"8��e#���r�X��7���3��l�a���>�����s�AwRr��t��q??��}.�\i��ܛG8D�}��?�C�j�n���Ir�3��m�����귋�+�f��*]�D w"1d$����U�'p?��P��j�Jg�α�5��H��c��x=���"�ݞ�08�^;�p����v�}E�Z�Jt�K�V/�ra�3�s�@<�A�1�����[�%K���2�@.s%�+Պq���,$/���i�}�ȞE�?5~f!�^sa�׈�I��2�G���� IS�FW0W|1���_��NHM����6�`����)���o�����'YD����\���x�>��T��T�D��=+ۑ�i)9��^ٺ��D�p^c���e�Z�� ��9�KBl���b��l���zf��{��'@����o�}1s���a������s�:bu�<.��MB!�M��!3 �lz������"rb���Бs��ˮ�l�j�&P��_7HKNwIJ&]Zæ6�����_��L��gU��*��3�d�f�Ւ,�����W��+�.�g�	���ql'��4�����RX�3�.�z`�~�A4xk��{;�%� �{�����vB������V�{�g|j�.�����
�w+��9B��OE��/���V��!�_T�q�b�?��>#�ȉ9Yy��A_��͖�EK�Y���L�l�#H^�<I'2�Qt+=���򺺈�b�]�(GEy&0��z�ex����k�.�*`4�j��3�'�c���>����h�:(8%g$9g*�F�,�s��-����{�l�m)m"��x��M�9*5(�r�T1X�����S�{��0��8����D������g�ȭ:��� x��e��Z��0���@��>][�wh����ȴL���ؔ�c�G�	l�$�pTOD]WOk��Q�5�{�=�R�*n_/�6X�V}��"�����}��x�<�s7���_O�bg��E��+��$��	���k(TP��^%�Y�T��P�����y����e�oא;;e���(Z����~���
�8=Ӯz��P%�����Ɖ���!����N޿~Rb�<{�`j�?�k�.%b��f�����2V���7��O��"�p9��EkOo�:El��pN{�d_���G�.�'���rk�4�a�9�+�����Kb}�n���DÚ�:�C��"}��DȪ��S��O���o���>�쯥9@��ٶ�ހ������Zu��$!�m5/�ϐ��O20;���iɾ{ܣ$����G��lv�GrGeUy�6�J�P=�q�r������Hv7�<|J����n^��R��	1��K�ĖR��f�5��Y�=�e��'�x�E	��{ɷb+�o��H��I�TY����.����߈�\J���Y�b!��ҀOt4�����M́�s�ǹ��dw�r{����"�I�iչ����;>+�z��+8��eH�|�Qא�6<ᢑ�asx�����N�NuO�~�"_������)�ҧXL&��W�m&����	ϋ&5�Oq�C��j���.�w1�-��/=qX��}���6����~��e��ߟcW����' �n�sE� ���}�o?�o?�4z=�B.,��ƣ�Ӽ8c*��?-�?�B�����!F�xD{R�(EHZ8	��1�c�lz��{P�O�4�#������4���}x��т��?�s����Z�8�c�So���r/�0�wXW�Q�T��Ru��*i8n���{40Rk�x��_�*��U��_�]�K�:����LP��e�3��m2sɮ�:>
��S���8�H����͐�]#�`R@� �C���=�v��^��~��R
�>�������^
2�1�jv��Y���4�:?�XE+�/���`ȃ�מ(�����>�A�_ >9����z&$���>�%	��n:J��8dP������=��'��S]8띛{������oG8��- �D�4h����N��E�5��7��Ѝ�o��!ϙ��)�`���ڪ6�A��*��1/]�/	�
�~[�K|����N�$q�*XbG���4��C{5�)*��R�E~�W/��I��'�<� ٞ���0	ջ�m�����5P��Sg�)�Z%����o�:,�5%1�7X��9�q����/x�!��r��sw>�5� �@� ���z�Bdf R�[-A����X��ׁS0��%:�rg%]�����9���-��U������ "��Fq㈏�ذ\Ҩ��<bټ��sy= �3bI�pU���C�*]xy>�A]����?��w�15�P^��fWK��/ަ%�`tE��!r�Ԅ%?s|�t�H7�h�11�=,�H�� [m����/����L`T�"��uK����/��>�KZ.9E��Y���2�i�u��}��D�:�v�w�=2� u�p���E�\��PXY�w��}�x���v#��<�-����6~8��!��H` �EYJ��,�$�Q

��/�l�P��
)棨��<��$n��Cey1=�ZLX��V��ˇ��8�jNe}6�b�� �uO,���r'� �8�D�~�)���xT77������x�A	���t�e��4q��x�Z\��<pt���z�\�i�:���������k�#�o�U%�GN��K�7B\/��
`��?����=�8�h^O��?҄Q�9z=F�"#�g�Q���������z�x(���V��$�t�5��)��-�9H��4*5�Ց������SMm�Q-������X���z]w����������~]���z]���tZ.�M0��g�۫�� ����E"����Т�AġFպ�u��6��{��sH�]��F����+��p��L�<:r~m~>������䤢}�¬�����7#��;�e<V�>��hD���:�	r#���8Ht'�$��x��!�t������o�ʕOJH\��mE3�{{S&�ƍ��L�]҈�d����-hq�t��^��{�_�-7?,,�g�]�4$�VP(IwQS�[�+�>�]�k�nb)}���/~.&]�K& �/�l�f�~�r#c�^���@>Xr��it����g�4�3\��M'�xH��P����l�����_�1^~w����*�mF+{��\�@N.b���]5v����V@9�M����#
9�GR$����fD���a��4Ĝ��Gg�?��x�c^4r��%��@A&��a�i᠄�X]�88	�p�Lc�<Q��b	pi
��U�oe��������{y�OJw]D�C fk��zm�Z�>����A�]��}��g�:A1w��Ee����^6B��I�����8���ؿ*YZ����`����E�0Jg��L���J�'0-��ʭ
�-�n-����Ȭq�ԟm7k�cN��u�$�KQ�
W�j��|(+��*�nLw������cb���q��Qp
�3ޮ�Mӎ�ɩ��Fc����������`�S~w���m<~G�n0��,�B!/���ȔLː{\��Dt�q_�%���T7^�<�:Er�	v4����l�	eq~�ʇ�����K�D�,y�,�+[�"��YO�V>�|5�\��x���N�� Ρ�y��{�v�7�i���Ga���ܵVJ�/2��F��W��u�����&�� 
�9�����B}@J�G����!���O��Oz[�/�{���9��s��X��B#�p$�*�v�x�A(
�w֧9��I�������ޮ�Z�,H���<��]y�U!���_�ap�{��b�=�B��֞��a�aM�Z~��i��O����r��6R���E+��K/L�xkoQ{V�a�%b�k3���C���9��|�i�ŝ��Y�hX����N��W>�J���V�t���U���YQ��l��QW��vZx�˹����j�Q��D��)���6����S���vn���Lqbr��������k?��Me@��'Nm�'����R?�v}�_a�W�d��[n���:���	'=���=������U��^g��8�bU�8A�(�ȿ�0��.�WK�ޠWz�_\��v��>�YW�X"�Ѩ������L~�"�J��p-��)�d�"�!{Xc:\?s��yÐa����ǧ�6*>�5����qS-h�ڒ�B�,FW�e��������wc#.0>�<��o�W`jl,^{���%QkM?��vK�!?��H{�q����Tj�p�D�ݎ�{�M��2>��x۞f���&�ˎ����ՅNx�ۚD���$�d��IF��×|���q�R�T�Fc�{�D@cЁ��6�\�6VG��Y���q{VG�z��	s�c��h\E��r����v=�a������b?/�<t�]��-�$���g��POʝ1�ud��u\���+JGV!ҌG�O�����+��ri��z�A���&È�\he(J����Q�h8����1ΏͶ�8����W��6�!�֤�����E����im�UL��}�1Y�N�pk�~�d�ڔ�Oca3��Uh��o}��*&�ܴ��'r�Q�i{�|�ܨ���0 �G�qѕ�c���{C�Y�t���!&�Z"^k�
=�k�f����*F~*�&e3�8��D�y�d?���o��re�K���EeM;G�����,��Z�o���P�c�#h&	#�R~w4�OA� �\d��)��|ъ��+J���/uE��W�V�j�3j|I� �ױ�TL�t�i�����6��Lh��V7H�^���D�z�#a~�8O��RO�
��⅏k��],P$׭(��*ĸ�v�_Ǟe=sƑ'�\�S�>8��W�64���&�f�~�o���x�6`����~aW����o�	�r��"��p06�b��΁<6��N���Z�?�x�H ���籓tؽ�O�Kw��Vso��둗�Ak��3T�rL=h$��)����nN���m��w�����j7|�+�O��A�B���~zg�/����dJ�����BaK ��8����ӥ��	$�[_"LD��E�W!��ςcf��D�`-�i�UL���]OD���Y���9��m���\P����X�L������*�����=~�̙iCF�4�I��f���Z������:���G����Ao��U�ϫ�GMe�n"C�V7��G�_�
��PD��ƒ\�g
�pC�RqX
ڟ�hz�,��C;X8��y^��\��D��,)'YC[�Iw�����ze���S��[n政��u)��<TL?_,���2J!�z�y�� ���Ӗ.Ϻ�,�3��d�	�B��r]+.[�л/�mCB�������<���r|�L>���/��],����`=M_�.��ր������^?��ڹ�` �^2�>h&���q���P�x��g�T|�)vy>)��6$EUwU?�<8r��Ϲ��uف�����^�MYub��)Po��﷙N�o�AK����@��Ӫ�(���.l����%�/��,d���Ki��*�ǣ˙\��'�L2fY���*rҙ���T2�r���Q�t��M%5�+��H]P�Dk�'�ݽ�vJ��>���U'*WP�.����/�'�DL�Mj��)�z���w�]�d�0�X���Mqa`e�ߵ,6��w��MJ�����c����F��YW�S��E�?=��3����麌�Bk=�K�.+���wwe�UOπ�@�?��`M��Fv�4C�����^���o�����e�����6��%m)�E���d��⒔f��}L�ɍ���%	��UM�ؐ��y�y3�@ꒁoI�④r�UZ"��lAhr˔�x�]q@yD.h�@r����Яx�t�X��͏��������LL��N[W*����\he>������0�yd �!q*/9p�o`�����*ab�bBr�?V4Ϝ�M����37fZT�4̦�Ӄ�L��g�]�9��o@��)��zZ���\��R����w�y�h����v$A�x��<M%A���H�H_Wi�#<�z�n�Z��>�^ɸ�!X�'���o�jW�~}r���m��P�4-˛.͏`3��+��L��.]I��q�F��O�uІ˞]~�L�W�H�G�.&�g���Zr�zzeF�Q���ۄn�C���*�2?�<��g�Í����H�%)(�-�C�1�#��E�e8Vzd�^l�5lNo�G�J�26�h4���I԰E�
�lR�xq�Ir�^�Dnr������n�{5g/����SGn4�ZŽo[�_v÷.=8e�c��nu6�"��X���uA�A��"��f��EZze����~4yD#SoBn��wŝ#[��#�*��y�%��Hr�.A���f�\����W-Oו�`���@�9�5)@������(����~h���x�?�9<���'~�!���X�W��M��=Q~�*�=	�(�}�;)=�Y0Q!�?����~W��p�{ދ%�ֳgh�D�C�T9{��nF��Y�fZ��N�fǪX<���2��YC�=��Q̺��r�N���8�t��G�Ȫ,;�[��8�!;�QC���UO\Od�!�n��cAt5�7,���Rӂ��ZW_|�󯤴;��,l"�XiT�͝�Q��J�獮��Ωx��R�М�0"�{�F{�TŒ��qV;Y���hh��vs� ��q��N��E֔��3s�j�6��vz �٦H^�$ǆH�����W�>�X��$�����o!�W�wpQ����ug��K�ckrq��'�����zyO[��?L��r<9���7D;^�t=�5��n���d���lJ��OvͶE,���I�v�&2���U%LJK$-��I��������U��*l�/����篏k:"n ׿H�]�o�\��~e9�M�%hA
�攔��з�i�뷓b��A�qg��u	��awY���('ϔ��v�]�4��/�^C5��Yc=�ˍ��U�U��DC�5)-��B�**ý�h���O1�'�{�!c9��������,�c�)��yO@�Z�&���0�2����.�J4������NCi����Y� �-�^v��,�IvM�ӕ�c�ߐ�)�E�v�ʼ���2�'���Kʎ=�D�P6�mZ_&Z/LcK��6���vM���ZN��.�6ym��\��BV������o�}����;�ci�Ip��Y�n���+,�l��|	�z(��r��|&+������q�w�9�G>֖uس�̠�Y�)�ld��rM��Ӣ|��_��K�ݭ	#g�~�`��N�{��]������]-���{?��К�tK@�6�h�K�9O��U㲗SEO�y+!����z	J��q�R�h���O^C�d��&����c�5��M�?i�r��9�|�5?/�z6?��'�\פ(�ޏ���=�Z4�hqLJӌ;��#�Wu|<W��Co���`u!LpSy�y((u%~ԕ��Y)����" ���eM���r[\�3�B�2b��K�`��t[��`����.5����f����np�+һPD��ۧ�i+K�O�aI����!T�l�,M� h�fC�4_�S��4zWS��N�_C&a�G.o��߼$_��VwS�%��4",���0�c�LB����X�zl^Ŀ})��[�50I[���\�P���~����P&%®V|�)����;�.���;�X6Ò�n��=�����,�4n�U�O@��K�ܸf��C�h�/ٌE,�Q~l��2%��cG@����������x?�A�A�X����2��A��Wӟ����Cs�"?}���~�������H���D!��~�b���%��!u�h¬���؊�d�6�QG�v8��{��;r�d�巑��������썻�OKN^��B-���vUBv6�n���e[FD�eee��p�W���iM[aQ�-_�eQ�W�|Jb\YS���,e�?��.D��422�#��vy�$����k��^�2epy�(YƗ��-�%��\CB&�\��%�mc�;h��4�#��`2��1%���(�Df!��4tM�Y�ocW�n���|}+�U=zT��QP8����N��%,�Ϟ>�P�=Z�����ۗ��p[p���XDpx�Xz~�����΁-��>)��VU�[Uz��I:�~�GȻ�nO[1��M"c|@�"�R��疖��4vD�@�#ig����v�c�����a�E8��S'剸!�GC��MU�ZS�eK*5Ǻ�t�%��d�"0�0��3���*پ�.>]������iHK�Ӌ����u�T��!�k�!Q�j�=E��N2j�P.� 9����@�e��V�p�BL�ړ��

̚t m?�m����1Š��}>���6�.)��ǓǮ��k�y����K�R����D����0�ӛږߙښߙ[�%;VP�����7:���%���w��lVRh�ҹ��2�:qִfgZ�RYO6b�4��+���Xa[y�g��zDO׶��b���j�zudb�^("٢�����\U�;$�c�����y+�ZU���&zjs='|�𱫰K����
����;[���b�+'�������q������	Y���b�	M��??;���k����m=�+ѓ/��*�n���;n<���_�ӦD)..{��c1J��CI_P�Eq>�ۤg$]Z��l�zX�J뒉(A�7w�{Tc(����5&CH�6�m;��P.�#W�M5���/3KG��|�e�a4-���1�P�rZ��K�!���a�����'��"/@��Fr��;*e=�R%�����Ȫ�)J�sl�.�)�ƾ��h8]����k _r��8��yJӗ��W1���q�vR�Ga�5j����Au[I�yפw�q#���`�t:籆|��$�IŻ��|���sy��'���JK�:KL���ƙ��P%a��*H�=�4-�D�DJ�����ճa���5� ��5�Im�G��
�lQY�W�|Ϭ�i]����G���h<*�7����{4ȫ�,��[l��}7�0x������Y��4ׯ��p:��+~�pě��:Фc`�Ԡ�iP�������[�����z���f3~o;�V�$8Mao,��iA�D�ܦ6��Є���e4�ee�I_�%޽�pz?�磻�����K˫��m:�4���'-{)�!���1�H7Aط�R�0�LB�y�f�z7ɗ�rz�a�,$�����Y��=p�Mv��m��[58V�r9�N/_�h�ݸ�~Z�L���4ޓ/q4t����+����e��@�\�C�H>��t�w�AOJ�@� ���X�p|k���ɠ��jd���(J7��l�J.�u�y��	��F�X�� �%��ޞ��U��&O#DKx����V�m���:�O��
iق��,�mC�f�C]J�R	~��QoX�pB~l�$nxVx��Z�)ظ���j�1��c�E�-/���3L�t��q��=��j�������&RH�8�h �}�ʇZ����B5)���:#�/He��dG�&����*�H�X���g�($G���@��E��x�{u�U��8z�{�m�^�����p ������i_ٛ����A>uho�+��I�f��H�c�\Z�m/��%���c�@��~Cȋ̮Pp2�;k�����?x���8��c���
ߞ�ᆓ2ߺ��`����z3�/���+�2D?�����(.����7�=���Y�����^�L���m̶����k�z��_�,�{��g�*��9�X���Uk��޴���x+��D�l<9KJ���Ƽ� �2N^�X����՛���3���DZ)qg 棭�~��d�~V��ƻ��^�R��m�S'�Χd%�U��8�
O8V�NIk8�5]���s���W��\ݖ�I��(ga�
g�v�S<	�ϡ�\�YPꭩ�=�dΠ���r�3���+�m�P����TIҲt!����d��Ҥ�ƠKܳaY ��ǆ�ϑj�:�B�+|��]�ʲ/�F~�BW�	8�1{/-5����j�2]��`?��яyZ*�.�ń2,�_h\���������D�����[N)�lȮ��,���D�@R���ld��i'7���*�W���>��\���à�$u�	�y�#L֦��.�
��`C�L�y�\� c���ͥ�P�W?�FC>���C�"=�J�ٓ�s&�{���(�WR8#�h��O�aj�$��E�K�����`����U��y�a���涁>��8b6�n����0��fI}=��!][����VR��K`�{/ �G0����z���R?��DPg>���*���O�G8*�;��7XɠkWj����0��$s���?�[[�Υ��K�=Bw ��:����G��	�ߋn��J��(m��F���(Ě��l���.Ĥ�{��qM��nx�}$<�7m]����l��D�d<n�oT)_iڂB�cʡ>%�_0��,*���\HVZ�:�'u&��dL���2�������/k�/�p�dT�lJAQW��e��Ӟ����ot��6_��C�j`+|�P�U����C0p��,"�0����ND�P7;���Ko�7�qM:�㟽��y��fa��Jī#JQ��P�]M>b@>���S��xiR��}�t��,A����0#5�՜V�&[r��C޿׸%5��5o��� ���O��f�=��/�8�w��ۍ�Y��ġ,�
1��?�I��x� Q��&)����Ē�L�f�JE^�Fn2��l����i&��E�&?�g)����O�ڥ�|J��o�-�o��gV'Y�5�D��U������~�խP�\��t�X�.O(�G�%��u_�u��ڊ��y:���?S��{��a��Z3ra�ݍ�M��I+���8�K��˰�������� em�S�.�L�&�����,h�M ���޳�/��^���a��Ʉ;��"��[Nz^j����b/���������Di��>A�YDc�y�f��*WCSX�ZI��ɟc���5y:K������;��S�-�n6xe�	����<�%���7}�YL*��>��X�^�P�@�6�8$��t�*�D��CM������ c�HD���k2!�+)m�JW?͖����w��lM����\!�j5��=�RpI������r4��b�%���o�Fn��tZ m�5p��!��x5�e�Gd߹�E)`����=^Vm�B��pz+��5�3��Z� ��ca��O/ 09�;���I��ތ�O��z�&�W�Zq6%C�oGw��:��2YGpV֌k��F
��U�f�AM���m�(���?�^(�|z�W:�t����s�s���E.����7�#֖O�}P�wd�^Y�����,./11% ��Xv�I8���y�߷�"u��`ܘٯg���i��AI_=`�s�
&�&%6�H8�����ᑗf�V<��OOΈ�"����\Me��2�5�q�Z?�J:^�t�H���A �^�+(`��м�G(�&[���/?�ɊLj� Mbƽ�~4�mN��zs�@E8��5������66֫����_�5����( {�G��p�˕�U�U���ǡ��{77-#��u�\�r�������1	����=�~	�|:�k��PRUEg�,���|��g�^gc��Uw0�nt���:.[\��
����bCy�sZ#�\�>�^�i�!�:5A幮)��J������T��������ʲy�=�OĜ���z�"<ח3��r�JMgg1�6\v���pw%Т�=��U��S(VMn�����t��I�wњ6����1���I��Q٪�����~�^�n�Z#�jX�GD{����K��=�hO[�Yxs`�g���:����+��s�9z�	��.Ƕ"Rt%�{�C���J0��M;tEZ���P�A��թb����|e[P��ʠE(b]�i��\ýϻ���y�F�#^'g�QtT6�T��.׏+26 a{=�,ǒ�5���v�ᅵJ̺�Z�|Ü)DB��#
X�ӽ"t%��[j�#�m�G�G��q��5+O������F�:�{&`o����/�C;���Dd
::��R�A�ׯk�(Ĉ�#{��U~k�A>��T��Pdvapo�����
���x�������w���%��7���_|�����ƃ��Ë����3�L�������b5�fQWd��⡖�ɑ��//Gn�F�����_E����ª�/ő�>QڍF��"��ǯ_[,2�rUJC�/u�ӭR��ѭԼX�5��gC]ݨ���l��fm�fGz錖��ƻ^��
7�jkkg�ߡ��k�ϝ��Q�����_^lol���#����6Rh0�m�-�f��-���
1[�"#��S�;i+����9���胦��kH��x�!�-+�X�)~4|����mDͼ�(�<�-�x�J�PoA}������B��~�ʘ�ƈ�)�IvȬ��
�����Mm�I�o���E~
���?!Y��u��k�x��'��ʘ�O�b�7ҽ�j���B��i�
�٨~�IJ�VJGtכ1���EC>��� p��?�q�_��R�2�6����As�x&+d�Ӹ��W D�����k~R�뢤���2�Q�g�����'��XI��t�xv��Hjg~g�bL�a^m��T����:���������H�ېV�v��8Ո�=ţ��jE��X	81mܜ��5��]Q!�$U_I��כ��'Ȝ,�s���zZӸ��Mm�TV�[ٖ5��i�.Y�Ⲟ�∱C:�=���.���;�SD�(�j|��xz�Wh(��Z"��w��>���~��ŝcf���#V�^�h�d��qz�kZ�.����1$o����5ɱCqI����#y�L��#-w2�?��B���՚��/�^������gq���R�K��
T���t�N�z님&Oqz�ŀm(
�!�D7�C>���{�稙�����E�4A`�\�+�u����h�{&f"N~E�54��ڂ��V�ϟ@�"p�Ho(ώ��ZC^�w,�ı��^�_M��D]�^m�e=&(�b����T���q\�'4���Y�Q�ʥE/�m
����+�A@\�>��U�`��]`12�u7���y�y���/�����%Ɗ|�V�}�V���/?�Y���T�k%��`X^�U�n���v
�=��Fವ�t���w5W����D�qC]��
JY�t�Z�;�;	g��[����B
��m�?/(��K^B.���6��)��c��%�ؗ��k}mV�G�L_`�s9fL�MNcCʨ��ID�#\c���z��������6�?���,4~Z���T�,����1R�d�u�Lm�V��)���_Ojץt.T^|Z�z�W���]GQ���I��@e���gb�3�����`ڳ�]^�?o���g��,��>���'c�5� ���&P|��#��&ٛ3��Y��4�)��>����R��Y�2�#c�3Zv�S�
wӴ,�����ia��R�'�� ��5RL�5����'$(�79�c	e�1�G�Z�;jW����:T1YR�u:^S��xq�P�{,�q���Xeޟh���oG/�Vr`3�GZs	�獮9Bs7�u��\7^?��V=#0��.�R8ЇQ�xP��r��AXM��9졷R��� �\��(�C,�����E��=_q鷩ě=����ej�D�2���{oA{�-|o�}��=�|�s�_�X:��*����C1qu�[k)R�v���Hw�3����;)0�q�<��hM��K��
�5&�Ä�|��uwF��A�a	L�B�# ��Ɋ�Β[�ү��!��E�$D���� sw�w�dH.3d��x9�Yw�7�n���QY�Z�9m��= �������{�uJ�i.����e�03���)نP�� �R��|��8�H���	�iy�{�O<��0T���r�:+>��g�9��~VO�#���j2t�3�2Y�����@��Ѝ�`,Q(��d3J�v�!�L�RmTl,�bݕ�N������w��5�K��ẒR���/�إ�G�h��q�S*�H�����'X#���U>��e��0�#�"�E���}"j�G�ǅ"&���=��{�\d��l{��tZr�i�N�c�����9R(�F��m@
�L��8%j]�6RT�����|�<�莰�'��sD��\�*���{�fۻ��4������];�p��Ή�KL����x������ќݗP��t	�s��X��T�Nƭ#�hsO�^2zQ��rBf���g�6G�F��|
Lf�_����|h��ۼً��"�<������>�F�ai�|޳���i؅��8!4�2�Y�(;��y9�����ĬV���c[gC�O��uF��xG��A[�`��{|zo�L�,��h(�?�a������C��Q(\�zn_�k_؅����50�h�m�
�:F&��5_V1U����V� ���g:[�v�"�����FiYR+�{�J�~��j*a{�i���\��@X<��|̲���l��k��d�������f3P��.����%�5T���#�Ͱx�����1~�5��X��{e�_�����~Y���7�u�l� S�f�ف��8�n�CC��3��Q3�AS��5���X<�G�(5����2�]1��r �X�A?s��/���!�(O����7���]/ =�Ȩ3 �g@���&Ê/�P.�@����L'ܟq���9ձBu;�K"�����w���^�s�<U)��z�l�r��R���[������O��#�{�]�&�^V�Ǆ�����/z.��������.�I��=�+���R�+\oc�O|�3䏝�������_��Q��u{h�J`�{U�����x��rv� �տ��2?����M܋�0Z���u�y�9�����ٝ�48w-1��P!�M�?>�?�h*QsW�X.����x׳zm�`f�
g��xc]w�W��;4��uF��P��l���F���H�;0�u�R���K�*Z�8�P_�2p7����?z!k��a/��|����/�*���I[1��x�e�l&������Φ���|�<ͺ��B��5��Ƴ�E��������m$�ۗ��Q�����G�$�d���r�� ��S����נ�,8���^�IAe�eA%�Pn��maJ�<�Ƥ!��>��Jx9�ķO�L,mX�h��q����wX���=G��T�&*.h�[g���r%vR�pK���K�N^a@L��ݹx%qa���Ǧ��^�^�7rD�/ôgy����Y��NZE���I| k3C���z$:w�b�9B�-�'��l��?��d������7��~g���|i1��T�ҵA���{!o�Ǽ3���m9��Åwm����^��*��'"a���px��k���7_�-�3��a��ƫë��)��.M<�7�z6}�11����Dp[��W��aM�#�+�J�NH@N�%�&�
)=�/�Bܯ��.�r8����;�J�/�9�c����I�⿊[������[|���Y�S�<����J������A4���k=ü�O����jG�s�y�N����>��'��#PrQ��l"�pHd�2^���2T�9���{.�0��K�X��b���,^�����6�J?ieU�U�+��)�� �v_k
Ѹ���T�*��jn��C�M��g��wT�[1�IƄ�PЇYh�tMR�Wz����n�~]��,�������$aK/9�Qfsh�P�$'5�Zjs���I�����l
��<K=j�"�I��j��^4�^N�'�IK�fͥ�m^���lQ8~�]����K3�<ӧ��/Z���ܲ��0��c��
�	:�ZW�M���{�$���zmcf[|����Gr$��<)����Orz�9�|��vwَ��stZ�~E��wt �0�!%���hAi�^a���4b��O�h����m����4n�hY��W��&Oپ)T*����kX��[?d�S�����J������UdDٹ���p_�"��[�W�1�+��%��-	.*�ώ����A���0�P���n��D߫������Z�#�����GF�7<Ț�l9�'pP�t%ɜ�7��lə�����V��A�F4U#i�6`, ����]!��g�rw�B�&��^#ZGL����j�_���ׯ�f�/���f΄?�9�<>��0�5�P�ey�)"���#��#�#�m��_{����4�@��љ�Waˊ�d�Ee�pgA׸-��]�2�����N�!�7ލ7᜔�Z=�7	�nM]ITӴ,*'Be��%*���<zY��YH���_��d�P�JM,7��30"�"���"�Zq�ߠ���1XP6�_=q�zҷP`j�M���c���(��r��ğ��ii.�U���_�0�����%{�c�j������"YgA�渦�l�=���x*!6��6��1��þJ��&��!���ٰ�{4�/�������N|���$�xu.�k㛈1�Ä�5i��R����~�<^^�Ug����H�\c����9��i�U�Ec4n���i��
�41��� ����!����TY��B�׳����K����)��!��w��T�5.�)$��d����1�S6q�7Ux?�m�<]��?��,�plp�j����5����%�.ׯkKhcT�s]�	Ǉ�R�NfJ���( �6�G��5�G��U���E��ض-WQ��mꆣ�%|�H�����?�X�����#U������A���-*(�56DN�.�H�7M'����'����x ��W�C���ׯ����D��
�$���S��`I�f@=leW��7l��0�j\�|c��s�_i\�~E��M����OL��������� �©�}ʞ��H�?��u.İNP���M�n�R_�r~�7|�zŉ SxE?�蔥T�t�eZ�y$W�����>G$�J"[�(Bx'>V3JR.�C]j�;v��&����NzpJ�4H+���<n����A�Vh��4R�\�'��^o$ ��gr�ޛZ?� �[��$�l�@�)��/���s9U�$���w�뾆�[#
*�.�z���d��t�4������*�g�@$gnῒ_�g[����P�\F�f�'�fD�`J����uM��	��v��1�;<�nb�Ƈyd6o/�+Ҩ�7��.�c^.ڰ��1�h�M�py�� ��4LNk5�a��[$ܦ��P�o�a�>���Y�+���L �����&����|�3�Ug����Mp�D�Z��N�l�e��V�>��\�W\�����a����9)6�RXDy�ti{����� ���X���L8·1��~4~�:�����Ƿ����A[c�!�]A^��5y^�����f2��c8fŴ7Fy�ba�N�=��	�j�#����[�����{�T،t��32?;n�Z+�r���Z��%�A�!W� I�}�W�+9kg{�^��T����o,
K�xH�ӞaupI�cE��xS�q�mU��y��F��/	u����5�rM��5���A?/���֣8>�eʑ�P]�Z��%��#����Jw!ĸu�����5�����jROƪ��]���	�\&~ GZ����[B%A��g��a�H�J!�������U K�������E3��M��@4�����v>�K��ohÜĺ`��j�'��c�B�E�w5�1��	�7����n�i�a#v�/䰺�݀��W�a\�N=��.`�V�U�LJ�E�ͥ���m%[��g ��xU�=�U.�ʟ�?�݂�w�e��I�Y��� �`�t�9$�A�¹l���PsP:�+����'�Z��5�t�Y?7g��d�|��g&ǯ���� �?��%�=N�bC8�}H�Y�{p����$`��#I8�	��0	'����{1	����l a��iL�,���4 a���O���}�w:��1	�tW;`���>h���i�.*���o�e/MK8-"�4
@���=|����o�g��M�UAEs���tq��g�Z�
����x�ʅp|K\�L�»���&������R���Xp�f���,|���Y��h��<������x:�~�]a���#�V�� �����S�flϿ�f����&̥���Գ-F��b	�?3�����(�%㔰�}�U�<�n��G2e�~�ٵ�εm�!(x�һ�N��$,o,J�}S��=���S���|�����y�F��RCa��X�14r�f���5��*h�-���8��� �з��a���:��/<���?��OK�OS��$��Z{+A���7��(ȯ����v� �}�!;���ˢdP}��%�|�4hY�b�Q�O���)��2%غ��%c#Z!2b?����:�뚽�Q<_]�A+�G6.윶'z���t���ސ0�Ϭ�4s]�"p�t^�w��=����١�|�c{�[�omڒ���ၡI�2���'�ٍ_�H��G����ҝ���_P
Rӷ�sD^4���}dl�l�#�����8I���Q�矐�t�}��<��+�S�?w��B}P��w�d�x_sP>�>o��9�qכ��Π�XJ7X>��>]}�O�N[_q�x;�uG/�Z�k�d��x����M)i{n��wm.\NU�S�����(��)�(a�?.��l�z�o�ɾ99��<p�իz�P��P�z��Ñ�}�P��4fdLqjzB�̠k|��H�SjwQ�t1v)��1Fk�L���?|z�5�j�aC��+��
X�l6<y���C�K�\���;�G�B���캿@��um�\p�{fS�:Z-%W't�/�����S�"UI��$,�F��N�l[I���![Q���Q���Kn������Q��Ypx�F#Рʹ�!�����<r}u:�_��&�/?P@��rgc/"��������0VSK ���<��z�F�/��c��B͵����O�A�:��9 n�����b���s	��va�~h #���m��3���8��&6f�\�I��M���Io���v|��ኊ��q�v�M��� ���L�� �x��~	�c�n����П�#m�͐%����{�c,R7N��{`��p�:)1�d�v���,mp߁'��	�;� HbE">I2��`{:N������4��l�ף��-!:Q�쳓����T��2�5k8u�����j	�3��7t]&�Ґ��B�o[X����xqU�!�3��M�|��OXd)�~E{c�s���e����Y@��-� 
>�!�Ĕ�oJ別^i3j&��x�"(d'`\(�R��}��l`��7�x�? @���<��4B��<�j1
.��!�Lt�y<?;�%����W�zr��e��5�w��W�~�p6�IGR]�.q���*Չ�%��Fy#௒$�Ulۈj��7�����?��ULka)$�VB߫�?�=$�JN�c�803t>%�7���L|��i�I�͡� ����d�,�o@}8�A��� �u��.�Ô�5�i�5\_���_䡊!_�q��| �ngL���	ݾ���͠x�%���6}�f�m���G �����Ed��B�_�m4�Y�L`�{������A�HmȌ������Kg��1�2�����,��;����`C�c(>��
f�C�t��-�F��Sא[`[T�
����� ik�PT��F���̣���s�b+qf��'�������|Cv��M"�y!8d-�����#�gC�U������_ �}u-@�%5�A�����I/Ĕ�C�|9��Sߝ�c"~��qo%[��a|���Q4�o��F�+ޜvZ@���:�WVa����6�GU�l���.ᵱ1���,,/�S���?j����	�b��Z�!�T��e~��0��R	�GwNb'��r���*�I�0��M5���VQIik]��-D���p��ڎ	�!Im�~��ʝ�&��Hu.��ؘC�$j9
�2U\)�*95}���&��o$��{+Y�W�9�,�%2�`r�L㚛 $U�
p�"R>}��Q�(�ߋ&�k�����Æ�C�K������>�D��*dX�Z��s�O�q�����;���rJ��m�p]{�$���΃"a�*�z�cg��D��!��:H���t�P��M5%�D ��L
^�#\e��ѽ�R3x.LGGA���U�p�Y�[+����K����!�Ά
	H�qc58@H�sLk�h�w�,t7㾟T-k��w������%$�ZwA�/ӗNK�{�i��щÌ��$i��>���)��w�:��=oSs{,�£_)�/���Γ��*��k! �E�T� 6�����T�&r�`I���˛�# ��ըI�"�~Qw�,|���t�C
@_C��:��|(��V�`�8�f�`O��`�?�G@/�0ƥآ�X}�|F?vj=����^�t�����~xv��j��1P1"�ӱs(�C[��W��m�_�QNH>w!Gp5ӵ$D�/bB��?�!�|n�T��RF�d�+��7(v�w�6YX����{>0����7:����c=hTP8�^����F��N�m�H$�D4���܇�2���66�߯�+o�����͋�')�Je"@v�L4��p>�����:T�6s��.]=HV;ޕ��*	6��I�c'�e�$�8N&~�A'�=��u3b,D��pb�dY��O(�J��"'¥б��wv�����/��!�1!����K���`�*������BC�;;;��8�02���L��B���1Q��@.'��MMVL�i�*eHs�;e�z�oX(���w�-)V��`�oÝSq�S�^��:�p�X��Ռ��-'�e�溛��l�r�x|��=��p���G��{ͭ��I��|lCCG�0 h%�>8�K��e�]\�͏���ү([�*������7�e�w�Ĥ�öJO���%���d�*2H�Ȃ  5�Q��Фu�5��2)��c��К����Wf�1*����nA�YapJ��ئ���ɽ����&j�ͽ&dЩ��p��I;��I\VU�3r�a��J�&�3�I������w����Ӟ��Ƀ�4�E��yap�L9�m�;��A[���$�8V��˛�*��5�!,�)�X��&�VP�g��>�ӗhܛI{��;a�rP��� ���2�2�EnK��O
����/���x�d	�#P�S~ą���k�D���?���do*�|Sƛ��'�	���
iw�u&I��
�ѧ��*5��M�����a�ȷWVvkSa�"�O������2J�gk����B����˯�.�oe�h��[}��٧�.��<������ kD~)��
�����g�`�5	Xtrg��7��������?�*���6�����ԍ���>�VUA��"���K�R��r�Ip�ߛ���mѶ
�8��bqt��D3� 	���4Ữ�-�
�z�Y�%^#�v�9�sj�f���%km�P1Sˢ2K

�N�0�"�9씷.Gc�P\�-Ѹ�d��"��i͞=�i�d`~Ӂ!���e!�٤{��aw�2��� ��N��=�O
A�1h;��#LS�����\p������(ԝ���g�M�v��z���N%	�뢤 ��~"���:\�&��ը�5I�1DX��q/��%�����K0��|/hmb�~6W͹{��{���p�,�H���q�ٕR�w�K�OA�xB%g����R�>M��(pȃ�R�B�K)�g�����{���'M�ei�M�A/B�f<J�<J��m�]>b#pZ�!#����ܷ�%��"���@�4����U9����0���P^		��s|��^\���������ߥn��F���b,���� ����d+�{o��"Xl�BoQ���h@ZP����� �pff|���=�ع��5k�S�3��3�'4m�If߹�}<@"�~>ww�00�1�rO���S��>=^��9���D ������
d����Ԫ�C���3w~����|e�*r�1���9``x��mFg�\�iA�n��)��&�\�ڟ}�-���v�M�N���b�Ц�{��-Ӡ���-I]�(���y�o�1Cܵ�qy:uǤS9Jr�!��C*ŧ��.dȚ�����a_3����2�� ]��*�����h3�lS�`�`�Q��sNLB��$��z#�~�s6q�a+Z����� $ei����*3hGV	B9RNHJ�Cw8���^Ȝ�� �w�u@��j��&M��ѳ���pG"�����ϥ͚�Y4:��p�o�J�E:�rY�4<�$��ݹy?� 2�*2i�[�e�$q��J�$w��[�\dͅ2��f|%�)���H|�,��추��}�9��ս�NJy	�=��:V�9@�&chϕ�EL-Rb ��Ms$B�˙?��P&}��P|-�j� @v� �H��M��7�d!
x�Y�S&L2)�I�r���hpb���{a�I��|��Y�k�^��
��ۻ�%\��j�<�!x�ߩ��'�[P�?ޢ���9����Ѱԁ�{�4jPٿH�.�S��I�%��]t�"`�i��;�6�>��g �[���ʢ|G�fAp��ئ�u�tA�2I�:�PJ���3�,��͆��1���#0f���~��*�X��G �v��c�z(<�C9�&O`	�?ׂ��=d�ٺ����F����r(h{[��Hԃ �zx;\��)ʺ��o��n�M�k:?@�!�c%dո�
&��M��6Gʹ^�Ƕ�c�m�?�i݄&<�N��'R�_k�_�@�:~�����QA��{BeF�t�e|��̤}.m���5����ʡ���c�n��T��^�?��ѐ3���"6��7i���̃��5�?U�C3h�-5ݗs;����̆D-�r��ѭ�S�_$�aTpD�c�63��N	���WZb�zG�!�r�#����.�#�{+'�&���Ğ��A���׼9��G���'ό���T�Hh�Y�U���n����Bv�ԔJ�r�����Ԍ;g�>��3���?��jI����Aj�b�T)���,{�fr�?U�Q�0�*_i���9}?S�[��n�3�evU5�29�� {M�qH�l��F�ѩ��pn���n�=pJ�#��2���/{�ހ�ɟ�-��&�X�@�(;�C��D�&�Ѻ�nkT|����Gݧ���ly ���՛��U�
ۇ�l=
S�S�,lqm���wA�Tp��i����j���'��rP4� 9s��M�� �k|�U#J���]BB:��$��,Z�?�]r�E�JI���Ͳ1���&��>�����B�D�Af�G$ M@"ܴ��&l�b����=h3:����p�w�B����x�x��92@��� ��9~�i ��T�\E�l©��[��kιr�T����V������ߎ�;mm�eY �z����`�_��N��9,<��lتt��1�zjzň�|(��\���.;�(�*���4�d)��g��z����o�f��u8�J@(V��������{`XA��"�gz��B�&p��:�F���V�[߉e�:=�����%OO���3�>�at�ڳ���>��]Pꘈ���,E�1}�P~��5��SK
�}�p�8���v�n-􀱻�7!=V��ͶJ���VZs�6�F�kF��'J��)�@7�� ����ݦsy��ׂ3}{����n�9�������U�vg7�k�< �j���Í-�`\RӀ��;��a�u^')��NB$"�K���*]B� g��4Gd(��d�������M�4��[m�e����+4�7�-��L5)�:-O웂����p�''Ѐ�C$�M�����p'�0����r�?޷�����Z�AR�� �
H$��!���̜n�_uғ
�|�S�zO���1����n���ڂhԡF�^t���Ϧ����Up�t��g&X�� K(��zE)� ��alV�I����d�\��j��$��V� Z؎󎎏�?�x�05���fWj�#����O�_Mڋ�� Q��R��~3y[)���ځ�յ��@���ho����_<r����Dp�MS�oɝ51��xÖ�:�J�Ts�����`/���t�Ml����p������
��{��2e��R� 
�~E8�ƅ��i�v2��kh�Y�`�'��#�z]"`��$�N�n��u�M0���5J>$���� 9���0.��P%����K��Y��T5�g� x����"V��)������6m��n�X�z�\�@
%dWzŗK�m���L�k�T<�@����5U�z��:�*��+��c�Sf���k�������PdM����(�cǇ:Du�x�_ �_<"�<A��^���m��"7D�t�.��9ǭ� ��e�fQ[�^]Ȼ߫*r>U��%�d�iԣ�?P]y�Al�5����(����-#����}&t1 `/U<�1���C�|�qK�b��VX%�U��5��ѕ6ˢh3Rf�
��2��z)�zD˄�����P�<x��E2D��f��7FZ�c�Љ�#T�J��vi��f���������	���y�=��Qv�@r #�qFqS4����͜�4��$w ׸|��N��h75H���:�GI�8[Tv��p�g
�_�Ƹ�Tp x	�c��h�y�dǥ�*��L7��µ��=Оg�C[2[�~�����7`) ��Wp3�c=ɕ)��%��z�+ '�x�����8���D�.5܀�W�y�6��W����֔��O���S����R_�Kؙn�ưJ��%Ĝ�20�d���H�b8}�%gu��5b�"PD��'���O桡������w�*�qʶ?ÚV�RX��H�E��kof'�SR���<ԥ�<�[ y��&�W̝��>ʥ9]6�~�Nٞ�r?��WJ����aZcO�ng.M�F��֤�J2�RM�����qCV��F���c?��WOq�c�Z�e��<��s��]�3��ܮ�:�+Uc��1EӀ::�?&z����b!M�Y�C�$z{����̨wΙ�WZ��qu(�������l�5�]���3�c<<{��Hcy2�����sg8�~&AKъC��C?��E���ࡖ���ZL �D�R�F����C.wzY\T=雵�O�l�!u�
��e�~��伳�� {Ƿ@�O�G&ږ�V1:qfʵ�D�Oq����g��^�h�̭��f����+[�f��X�� �C��n*��ѝ�-�6�U�%��!E$g[ߧ��p�`�SC-�~�-���ț_X/_�tx��D�x��b���z�´_���3�I";q�q����R�_�tpeggP@;H����g�֫ �N�4�������(�t�D��X=����zH-��Ъ�&��~Ѓ�����2����s������1H^05rͻ��0�^
}��.�~ƌ�%v�V���EhsK߳��s�xӕ!K�I�Piϱ���E?E�AGX�#W�Ҳ������!Ẹyv��UX��'�#I�qe�ރ ��J#�$˽;�4n=B�M�f�W�xޱ��S���.���� IM󰤣Ϋޕ�wLf��+����� uȕ���r�d֭ȟ����^ P\�#���e)�mR�AySa�7t�H�A�L�-�Xي��bE��x�  �	e��=f�z R���	ߋ}��#�$�[ ݴ}�b��1�|t'$�m�W}c�uXl���>������i��j�[?�Z�X���X�������&Lac�g��Ķ��u�a���|<5m[㍼x���E�afoȱYw٠V;a� �?�]�^�8J!I�pTpa <o�+� m��do��:�P���Rt� v�E<E;q���Qх~& ��e��1�DH�y���X�!#�{+izA�u{��mk�c��#T��R&���$Y'���P�J4�k�rU����E�Z� �x+�=��5%AW!�_�q�4t�r=$�Y���t��5�(�y(n}	꭭�SfZ��6�ʚNhH��`�V^��}����`@��	<����> W?�:����J��{Yotjs����b68:��p�R��+鼖���FD�z�:�?�J�>�q`P��m�0��-ߋ�~�X��w�$^�L������$wk���$�T��y�7n�ܠ��g�Fj��s�T��`�� (U���_��4;����#3�,���Q�u	���q��3��sO~'�u؟���)�'�i-�N��a�� '�ޅAW��@ilb�>��8ٵ�T˱��t.��<����]�m�0��>�I�M|��W�5�S@t F�R�)
���Vg��y1�:enq��Q.[��Y�P0ǟ�AY�6U�i�@�J����9�
� @<�ޥm)����A$��^��5�G�K犯w�f��ʐ�@�&�H`�-�{R��ޞt�,0Y�� W �Lo�C�?�Am�i������l��+�y���JP��nj,4xZ���q\G�^j4!���H� �73�6P�UO�����
U�>@!ͱWa �JL@���q+�_6d|�x�g`!���c,#b��0F���^�d5�p��l`��̓�0��\W`1aWQi�\-E�Xc�ҟ�KΦ6��E��
��H�#nNR6	`���#4o�}�(�N��|'��ٶ�d-:B}54~\�Pn�g�V��\-	?u��˭���J��=�-������f��U�-:4�lx)$WN�&�����Rƴ^d�6�6h1�/0�p�#�r@ImB�-ԩlmD�lI�����N�����۴���`ľ�F�bW (GC�B+y&"r�����-hN�=�� ����/�u�5�2{�3n>�r��rQf�W��&���
.4Y5n/��_|��&�^�
�N�K`�ȱ��_�]�N��?�
B��s��=ɭV���� ��(�f^p2���}ǍS�
��T��ؔ�<�kX�5�;L����I�_^�.���y�ܑd~�Pc��y�11k7��7�:R��A�B�ˮ O�ݙ41���#��p.m3Y�P�R:W�[&S�>>�jS0 ��h�}�݁{~/k�%�h@�S��r�B,)�;j�ښH�� �_�N{�4�S#�R!��F�}��d�P�������vД��2�Ew滲-��.l��9���9p
jЂw>�8�E[��r�5�K��Vg�vOy�v6�J�,���X�+��:�V�����ͧB�(�A=�ߊ<�V�h{}�J�����zw&�Ԩ�-R��IS��Ky#��@m���M����C.�מ8���b8�V%� .0��]�%*4ot�K��N���p��Y�E��z��EL��yG'�ۣs����J	�͖��K�͚	�9�()����f���
����7�����潣n*�sx^�D����S�q�_���|p����������C���b�c����Zh����kZ�/������;j`�5�Τ���/́�:'���\�T�naCݨ������]���݀��Ш� ��4m!��)��J�?�q��1Xt���۝�7|�R)+N��|��.k��w���uahk}�8 ��o��H�5u  �s%���d�n��3��qe`��s�;����	g��{�'��!p��f�|2���,�F�}��ӄ"?�b/��9��u�?��xF�x|�۩�\����k]Ŕ��#�'/.tJ9���o�w�m_��:+*�Z�ڨj��w3nJ�
�����ް��>s�ӹi�Qs]#t>�֡h�V~V�Ύ����J�C3���,�P�5Vc��ۻ�B�+;�K�nwh�Z MK�+a9�ղ�Tܘ��{�~�����ߧ�T�;���-�m���&1R 1�Еo*4^�¼;!���x���-�>[K�B�#���L֢���[uO�3�?��~O+�\R��,&4�� ��ky���t�=��h}��}晊�ɞ�R�*��RE]�2�:�x���4�
ͭ�k�x����v3\����U�+�GTH��_VO%�~�-
ֱL/^^1{�d^���T%�˥�|��
�ZYh�\�<?�1^��c�E�D�C�Y�P�5��/Ȱ��(�}��TSJ�%P�=s�Ȭ�>C?���_(9D��>ܩ��#��a�Xލ-#��:��d���F���E�M�(.UѺ2�#�`�R{�t���u%����j�]	LS�B]z���-�Mp���~����k i�'�(�>�ixW��%�y߸Ew��;��X�߫������3��"a_����d �r��!��?i"�r���PA˭�$�X��4Q/4|a�n>�p�O��z( f|M	��#+z������X���z� �u��8`�!z��|ʞ:6��K��l^X���Xh�n�gi�_��I�GR�0��{u�!uCϱN���tV	Z/��-��.�o`�B�E����U���ec1r�ҞW�?_E�>7��� ��F�l�vF�=Վ�F���9�B�����	6���}fĞ�%L�򴒆�jϑP�ę���ޏ����� ����Xd�rV�404t)O��dӜ�è{��%�ʍ'_X���t����؉2[v7�o�U�F�aX/>��:n��:�2�y�9�.���5�;�<5o*�ӕ"��S�)��Дq͙D�tw��R(GS�����$��8%*�!����^G�ɾ�
��6����9�6��{�5��`��w��T�4$Ò�9��_$\�i63+�V���A�v�-K�>o�������T�\ڻI�@o��&�B�gW��V���+3�a�W�l�WQ�/�.�ڦj��X�)�%��6�����ܖ�ә�m+ʾ����xXQʣh,掊_`�KI�c��̱�Z3�~v}ʴ��O�����=�Ŭ�[ؑ���譄֌���^���SZ�������<+���	����og�����1����Jy/�^6�R�o�j���`��n�s;���{z[(ә,wzZ,G�c�(�=�YJ
�k��zph���T������N�ZD�m�\�ӱ`u�b',�����K��%�$�,F�w/𸴵�-�f>���WS��>6`+Z#\3����J��I����am7��K⼣��^�k)�pF���G��`t%���d*z՗W�!(�,��N-g�+��e�L�ٜB��9ᛸL�Vie��-�&z�����f��ѓ ��LU�N��bh�T�Y�k핲���+C�U��0?�'�!r<pW�c"P
-��Ni��Ḝ�����%`ŝzt%���H��2nhz���d��Ħ��QИbpSG����3�q��v՞�����\��.�T0+GKcb&��pw�S�N:U6���x��2V�0�^�A��h�Y(	|G�$& ��5�`ҦSH�	�#�	1��E�)�L ���X�E�������>s%��h�<,�Q�������V�>*�y[�ל��&��~4�ՠ����g�q���ϕ(o5$�Rb`�׃XЖ�4<�0�ٰ���4��@�T�I��Ř�eq�>g͝_�:?��k�9|�.-m�9����.�1�R��í\ѽD��z�L0G2z[шo1}IA�����,O�T �*�}RñFQ�M�������F�Wriʩ��ǝ��݈�P��̝�LA@k�SE��i�G{�aakj<�ê�h���S���`���)VS3}�R󰾺�1^���� '��j��7�bMx$
���c����oڰ�B[�U��Y�~�$TO���:
=��Ҝb�'�oT9g�g�Z��GD�q�7"�I%�Y���l9H$���+�]+B鲥�gjx���6ԙ�*�.����|r>�(�V'f��T��R�ĺi-d�,p��feP�wI��l�"��@��yV�m�yS�Ȱ�s?PRHܛ��kg]o� VIe�jl�)1�J]6}V|)��,<DŃ�&�h4�C�:�h
GK �:@g	<Iў���F��xj<�3���K#�7)Ӵ�	Y��O/<"�x�am�v��e��Q,�Xp���S�.�9�������%Z�Q��"B�r��sx���*�t�!�:%�)Psgx��A_�����^n������J0����7�W̣,B�W����̝[�/���/P<�+�	H��������u^�y��Jg�Ȋ�;}q%߫D�܁V(�TN$��z�\�{Lx.98���]�=|����C���2"��$�"TiI��Gj3]R����H��:)����%O���u����ѝ)�f���#Ո���\�p6r�2<!
i�d�������i�@z!����bzw��y���X�oXt�lCE�.C�Ԙ�Ĵ�t�e�w��ѝ����PTL�I�[Q��ьt 1�g�yF���ˉ�h��>/�N�2�*k��C*��Z+���C�OOȫP_m�?��B�rW�(Ժ^ײz���F�����r:�*��]��ϩ�	�'`�_������[]f�E��w��vv�U�R#ǻ,kiǰuM�
�an�D�+F�S��<)�]6�����#e{-D!5�i��Z�E���b(ӽN�����.�_�\�,w��Vr�o�� Żb�[��3m��H���`��Z������u:1?-���%�������qF;�nM��yg��2�c܁��m:	�d��__�P�^m2��4�L�2����x�]�^���+�v��^�� �@$�k��2��@U$o`��˘�	K��O�֐�s�Q�W�Va�.x��<}^6���@jG�x�N��x����A'��KM��"�VF!�e��|���f\u��.��(�K^6.��c��x�J=).6�1
�x�z��,p>�<m4�dt��9��a�&"�n�od`99*�o�ݏ�Y��[<xhN�������9<6m���)�my�NH� )���c�y���Tnus��J$r��B��3��~T����I,0M
6pwM�`�˞AM��欥��N��^�s!�)��C��pZ!ڕ��1	�M�7@9�3��k�M�Ba�+e��i��9�-&���"(�=��˨6�N�lMQT�cs���#�iXk��QQ�8I_��d9w�80��?������Y˧�3�>�3,��4^Ԡ'r��Z�WFzr��|���q�F�O��Ou��n��1Za��N����\����cf���y�;|��d����v"B�~��ؘ�>�<Hg5��ի 5x���1:.�x�S�����l�a[��|S��/��[��hH�!X�
 7����A��Ӹ�.9>i�],ם�?m:�56�V�jaA�<��n#��S&(aS����}2$����Gw�1�{��^"�Vi�!�%��������H�A�Q6(u5��>���9B�}���:��l��̼�fyrD+}�ۑ���)ݚ_Y(-R��i^��ǹJ7��h���%�H�L�?��,=��|�.��ȱ�ez�$û�T�B0M�g�V}Vh%� !��qf��%jwǥ�r�[9���
��L*�Ŵ��������]K+l4/�D��_���dN��=��Rc�\����xV��Z�Ra��ߜ�.b�+��t�����[ݚ�^"�Q�Bކ���g�e�>��[��d4]Dk�)����X8��xv��o}`��^pϹgt��G�e�!ә��NgG؊��eI�ʝ$Z�qZ���k�7$kh;��(��m`	��\���8��H7��6d��	���rw�\���/��~�����6��>��9s���1pB��j�r3BW�;�bò���^���5��9�.�3U��!�����x�|���^���?�j�4*�I�8>�k��摚F֭c�����F���-*;�����j�s����7N�	�	�@,�M��Ŝ'C��η-F {|��иEk�I��Y\~Br�l,@~e?u�]�V��ٝ��3߹���Ic�kF�FD�z×�|���O[K��Q�X���t��s���[���1տ]�N�ki(�n�ւ��o����
��Ϝb�E)Ե�i&8�|�����}יͯ�����~4W���q�eow�憌z�ޢK�3_��񧨭R��<��l��V�!#���Q���R�U_�D�����5�0&;��=�<kG������l�e���p��΁F���<E�;~�SE�i���S�z�=�f����4?H(\���\�_�o����*��좬xڞJ��������{OH���Ɉ��	�e��|��	�͜5yZ��7m�?����'�E;��d�>AR�T�uqZ%-o�����M��/>qOa��%���V��W^�ҍx�k�(J��y�qˌ$#��k��R�L1���&���,�e�ٯG��T�4^}A�f:2��
h۪0��]3��m�c�����[���a��dT�Z��y�������^5�EUfr����'�J>���	�T�ڞ7F�ǆ#]ɲ;UB�F<����b����Z�nF�巐,����F|��?�����__��aҁ�R};Ƣn軆��t1��fDl*}����֟w���)Y�����{6:�;�Ȑ���w�1����c�z�?�_d9�d_�5�H���Ύ�N!������*M/d�LA�T��<JuxF�P�r�PQ��/'z��>�m.x��4���rՁ����[�eR6w��ʛMډ��;���w�7<��S�<�\\zJ�&{ǡO�������/�z} I����}��C�zшL��5+���}�<�F��m���P,l[�{헑�O�0���.�9�$�Sp��=�k?��Yoŝ �� EÅ��S��X�̀���͆'�6���ƌ�]�������Z7�����Y��ܦq��_�}�j�s��7��3����8�>���~�h��	=�,�CcU�}�O���+#Vp��8ա�MN�AW��k`׸��{*vXؠ�Zpv*Oi�߉�O)݈����@};'-z6<d�ڴ���
�o���r���ڭn������i�j��\�/���=׌�W[.A�d^(�E������[����ڣT���~�y���T0�O gI�h��-�KN?a�	�|A�Ghwk��M���N�7���l�P?P_�����#z�\?�Zf�NR�3���{����;hh�!�3����� {�Ks4��[X;������V����<y�$�w=u:L���̇�������A����~J�ޙ��糎�c_�,wj-+ls�c�=`��L�oKsi��"�x�ݻ�v�@d���F�3sv�B���S9J|Ď�E�5���,<!pE�\H�U1̥=����2��1��ma��Z����~¥!*�Jb�2�:�e����4�����a'�N��8et�K��K�p4�c�@Z�l�����~�*����3�tF:����"Q�_����}'�������~:9�P�=��D����d�O�M��C֥�vZ,�\���|r��Mn�ڙ�!	�z��󒇁r92Ux�1n�m�8_t������ʹ�@	��d�'�;P���2/r
�/�EE��~X�Y���m�8�g�`X7�c|���_ڤ֩���$�H�aа{j�����F�4_�NG
���]g��e�wq��8^�C�]���4��i:T05)U��U��O��=��H%4��t�!����S�Cή�sU_�܈� �a�w�kc5OE�ʹ�<�%���
�����}�z���z/(u�Q�گ��^�חp�ԏ-M�p~������J���x�����]��w�'+%�U�0�?�jU3s���CQ�h�g�&��̎L�J�bS����@Ce����Ye�E��F��G��U����1L�Ѷi@�^��p��������o��3�h 8�zȓ��oވgtT+#���v��@����+��A��i��3_�@�Q(�v����Ѫ1�����W\:��Q�Uo�9��v�W�U����K��rVł���t�tW;�՞�ʝD4ML�A9��J��s)��%w�Â~p�̝�3}Y��ހ�EY����wG��~���,���3��	��v��i�D��GN��B��!��U>��od��[���	�����m���6��~����h����Te5.j�9��XP���G��U���Р.�6����5p">�� a|��-F�1���s*Ӡ�YA��АW{U(��|i���'����?�'u*�
boaI������?�/A���{q�Q� 6��*uҿ���J0���4�2�riSşm�Mʾ�?tNuL��E1x>y�/��X�3�P�|>��?��K<̸>�m�r��a�<O?���$��M�D���l%���#�[F�)k�2g&���<�7:�p��u�Va<��� �	����&�tb��m
���m6���Óuv��Jq��� ��y��c
������!B��>@��I�H�ܖ��b<EmG]�i���^`�#��Ǐ���|3�DU�G�Te��s{�g������q�O�D�����]rmr��Hㆿ[T�ȁW�cQx4�;<����&�Ᲊ�!.��O{�\����ʸ�o}R��B������g0�;?�pR��K���aD����	*ǣF�l�E�e�������#�Ӫr���dP��e���ϱ�@��z��z�K����W2u�}`{�F£�6T�ڈ�ZU��GlR���̊�0���y��XH?��m*|��x�^�7�D�_�#�/���Ar��A�_���I�k�W����S��N	�[on�����?�ϒ�c��n(U_3�3r��M��̽�S�{jw��Q,�<9K3�M��ڞ�]����F�m�ork�x����{ӔX8	Eڤ��D�����z��0MJ�~����}���̽�U拆����S���N���V����{�,�%��{��G��'����Ny3$����R?��������a����X~GP��;R��s���J���!��kg�&5ǡw�<�`���o�v�'s���5���k�P�~� �;םS�>�0\�����DL��Up�/��Q��=����%���D����������˚���}.;��w�\�	ioЭ:��v�+�"1��`�\+;��|��m�D�f�gѷ'	ܢ���Z/�[ c�"t��c.��;���S�k��4<t�$y�1>G�%���Qr�{ȢylIz�-E�?G	���k���(g���Eh�TC��/GP�l�3��P{9��9������>�e��ƿ�:�����'����O�$چs#�ی})�%���Lf�$>���03<�v��mK��>��>GU�(��Ak�ڧ��O��X8�D��!m�l���1z��:�H9�-L����0x�w�o�qG$�*:�Z_�x�7�K�J���t/\��B���wi�&]�$����pu�
���s	DHY���R��d$�[F�j˛�0�x�F<���7W$�ä|�X0�͂m�ˏ��qG̻���iE8}�����`����9o�q��3_�|(U�*�օ�(3�Mn���"��g�V�֤A�$�ݨn�v�穅�9�Z��g|ޜ�x��Vy����l�����ُ�d^�e��F�/8��J�n���l���'�0�3uv܂�Rm1eLW���>SQZO�4(9�;�ֿM���M����'�d򟐩��7��_'���+��.S����9�x�����sQ�.e橿���d�yJwI>�pXs��PC�aǫ���2����E+����$��J��㳫����Wv�Xt$ݡ������Z׮y��5<R�x�ɟC�WW�ܐ�Zƨ)İ�(k�k	Lu���Fi����p��d��ɠ������M(��]�#r�~SM��	L��E�y���
ZKi�A��9~z�}��;D! ɛ�{�����ޕ��.U�2�ԯ0ye����8\�,l^8[���1�{��"��J�/9��"��"�\'�m��&1L��9�<��
(G�q\��`E���s���P�:T�zx�W�+¬~{`6�A��4؟���qM.��5o@/E7١j-�T;[�&�q�-�Ak�͟�C����Ó91�`���c}�FP�Z�^m���4�v����d�iQI}�z���ÿ��C�!�y_��/�V]�/�=nJ�n���)=�؂�R�^��W�x�F9z��s�l?`�U_Ӡ�|��?�U:D� ��@��{����%g!<Q�A�����j2aT�!Zf̑��y1��6��25I��B|M��4Xfb��M�9�h{}J��t
}>���1X�	E�!��Ft"��Wx=����I;�U��jy�h�.�|�
���;k�;��5R׬�����.���v���������_�$�~�yf�J�^�S���5�W��Nf�S��/_/.+cNMM�4�h�����q��"�������e�k�[@��MS�Tn��I�*)*�|��,~r��+���_��si)x�Z[[+q@�U�E����wFc�C͉ol�T���ȅ/%�(r���87.))i���쌳h�o/������C�e�3K��щaFy@X�֪q;���џ�F���ˆ+Gw>�������fgei��q蠩l�pΔH&r�������B������A�v��I�A_��,&+#�aw�hq�t�y�=�9B�؂���������N��N(�{�ʘ������v���%�;���эV�u��q�<�m��4���2`;�f�x�䅠�)�[�Ȓ�J��KtOq�f�N��?:.��K�!��U?U`u��E�p�s5��Gˇ�.Ec��Ԥ�O����4��)W��(�+`Z�����i��V�U�C��vx@k��b�M#I�{L����!�A��h�l��:ʣC��5��[�=X�)&ٯ��A���1<v�����+x���Ge,w~ �F��Sf>����"�o[���jB�z�|V�|�����wHC�?�-�	.���+�����e�HђKz��?����w��d�R��zG �#mk"�v��'͛�.\GPA���#�?��v���sL���� u��թc�@//�w�!�b�n�#S�����u*��'�|�X5��+Z��;�^-�h1S��%��B`�.B�!�{�Fd7l��=�S"!. 0�1��/	�0��&ɑ�䬓+�WN���'p��|-6�+mT��WA��[����و�Έ���q�O%)�$�ڑ*&0�/�F ��h� �rLN\���U1~;b�y+M���wD�T���i��y����u��WP |���� �R�I�Nj1"��ыk���X�:SGt��{a0ó������OLZ,�iz��D_�O��'52�l���td"
x���������~����)��@���(:��#�D���B�����3�t( fF' !"핂Ҫ스Up��:5( �� ���q�v�oc�Q7'q8�T]r��	/p,q�!9J��hը����3F�w iP���D2��F��x�<D�),i�,�����՚�͎Et�M�԰0.>t�`�u��O����0�����/tP�6�o����ԩT�N�����-�.��hB��kt�вګp�7FI��ź� �����~��u�h�<�34T�B�������:�>׼���UG'�3�- �Y�F�����?N?y�D�����b�j`�V[5梌��A�K����ccJN�O�݊��mO?k��Zs�i�g�M~��v�G���DA��(T!�N�#:K>��8(�鮁�lk6{r4���#�4�J�|�=?�Z%߾]�-cZĠ	hߑLEZ�h[�AI��T��0�Ù���NM8�N&��nу�O��2Euy����uT�J�i�Sj٠�s� ��J�㥞��	�Ng�/�}K�n��)�99�W{⟓�M��ݯDl� U{��&~���Z� ��(���ǜK��?���o�e3�=1�<&r��jaKgEÜ�.�a�o����Pz�|h4r꧀���0go*ʺl'�F �ڋ8"x���k�o��*���z��� �p�9]V�f.1Ul�Q���^X�h������U�2����
vS?��U��5Y��eu(=&�o��g����TGB�T��6�_�)*!��
� �sٔ���������'y*G��Y�A���P"�@,��/�yD����J����q�$��+c�+%E�ȱ�hgr�4$R~�KS�����*��� ���Eʕ>��H�Ne�f�g}����r�ؘ��ġ�{�b���a.�վbXH^ X��)�#.�kXnL��e)@�.Fr�,��+�JɎ퓉�eA TوJ���d��	]2.����(��c>� ��1�܄�7P /xY�IT�U��=O��L�\���}���O諾�XYpUޔ��j���W��w����.B 8gg�N?9V���G�1�W7�~đ�s��	�%���b�~���OG=����V���+�h���9�<�^l�V^��1Έ0UL�x���5f��������O����5������χy�HH���7�b�X5N��<�:�YYu��i�������Y��jsǓ���}�!Y�3�.l�@xSP�?���g����9�ޕpw �,�(�Tj�V�+DSk,-@��х����D�<ԕ�lI_�$���dBJ`+��a|T�v_���t	T�_�n9OQ�5��=t�<�,x\j}
i��\����4��F`Z�Ӛ��â����x��sT�p�*��	Siv���$�]�v�G����X�Gp��^�w� e�9��q����w���Gv�ǟ���qM��|P��RR4��pJ��	y4"��s�(�2���1��	�Ikh�(�A��s���>��FH�_�g��������ѷ_42I�Dw�H��x0m�9�kK_��4�\���!���Sx�s�]\�}@�4��7W������6�����D`1|�����Q8�%�>8F�)wcr�hk����:n��M�tI�	3M�3�t{')�t�z��V�	3�[VM��̴y���)8���#a�G�i�6r'�}1Z-YhIv�4�}��a������'ێ��O�<�G�f�b�c�
�K����k��<8�����~E�����'��Ø!'/�w�4kq�Q\K{�ر�W��i��/��(=$̍W�Y��נ���1�$���?�!`޽av��w_܉�զhF�1b���O)�E�P��<^�(��͎���*�x����7C!u�c�ku}�$��_�r����
�Q�-��������2�#fk~���z��g{����^�0[}<�� �_zu��n��9&�Y�q엤�#�/l�}�4��/�G&^ׁ�4���}��vb�z�X�߿�\�l�2]I�T$��C�O�O(�����-��ᖍ�����A�-���m��=�ֽ��E��!A�W{׏G�v���)�O�����~��l�u�_<'��8�յ(5i�ْ��^��.R�Get��^;a!��p/BBs�;�9���'�>ۃ�m@�i)NDY�QwEb]^�W}�ŝ���-L�G5a�[��gy�����}Gb5����'1�x!���C�$���c�4���M.(����u��#ǗIᴮ�k�����	ۣ��C=��'�T+$@�h��l�?���DS���G�`����_�,"_�$�jձ��8&��q�%�Q��Ɲ@�H٤����ax�ջἂA��Y\�$ZL&��)����` ��Y�ɍ�V��>���^��Ͼ�>(�4���3,�
7�<vp��0v�yp��(E#��]�lBu����3�h�#	'�r��m|�}LԹ��P�ҫ����u	������+3όc�{P�� �������/�Q�$U¥�/2���|nd{'��ـ��BM��`��oI/5���^��֓6�$T
�=�r@t�Zh��tM)K�{��]�*wo�#+�@/&��I�нNu�?"dw�UP-Xhf�������;X����Ŭ3�B���q`���	��)f[���҄R-�����2D�U�-y�7�z��<����IQ-�u�rY�������|M�E���A�D�0�&Н����p!2�M�W�2��km��Z ;XK����"HC���|�n��ˤ^n��Y�n��I�jڥ�au����I�&����B`����N2�vZ�����������(��L�J���Ȭ�Z�T��{��=��G�ӄ�Õ�~��e��[@�K�0-6AU�l8s�쑪�'���:������j֎{�Bڰu%�����"�w �P�[ʅ̨�`!b����ӿ�r<�G|�;>��z��'��$��ًT�#jT�·��S�1[��k���Lf�O���\m��ғ�;��|&��5�^���l?��mA��wd�V�"�K�"���'����BY�HF#���]QW��h��z�s�bq"�Gt��h��R��z��V��IoQ�!6����Z"��|�=��Bt�y���ҁ0���������#�/��R�(���7�/{��hn�+�
�k�zB0�Bh�;�=�\<� �Y�/����Z��LJ�ƨ:%~xv[힨��]���«��8x#l?��gߘ�0N�KMr���u��_������ZԴ}-���N40R�_�`��o"�� �Z��3B��Oj��M��:�.��(:�E��]���2�>,�^�ޏ��T ��ċ?��!��Ȏk��Bc�ф./�J���r;�Q����|Gd�)���)�-l��4��xf{�)G��;H�@�9�BS��QL��� _)�?�����t�i�e��q�4<Q�Hy����?`�<<��gUP(<�NY��F�_B����|�y�J-y3�q�W�"�O2Ǔe��z
wn�B�Tgc�e�q*���u&���7��!x��'"�c?�e����ۈ9܂-����6��u�^Q:�q]cl��+�B�.�f( �hW���_��ی���O��9Pe�[)���c
�}[/�Z��ӟD�B�p-�M}﬎@>�u��3��a�&�蝔�S��mxgn�y�m�%dE�7����-�ޯF����8�s��׏��o�K�V� gs�-w�p�'C�8?}�<��o��_ș���D<rI���o~㵎��h� n�z��-w7sӨ^�{yb��9��}��$�˘O^���F�J�#�ɂ�E�4��n�6�~�_ ���5ۿՀ:��(�,�C�M��c<>���]�
"!� ��4�½"1��C�9��-��{��+��Mn��˝�}�c�ps�L�U E�h!%ቚ��qɣ]���X�+BQ_)�C�����[�`��:00N{"�O^�dB;Wq�\���q<��Ë\�EZ���w���Wi� "�0N�R�0�&��wq!���2��� '�7঑��?k<��؄��9l#�e��a$,`�A��9���PZ]9;������ �O�R�<���,h=>{ ,<7x�  ���g��A��2y��m�T�w3~�0x9�0��l����ʸ�8��ݖ~���AO���\_]ഘ>�7���I�����P�o���!���di�ʮd�ZRI�ʖ}ɾ˾���P�.���}�$E�}b0��`��`��9��<�������+Μs��}]������>G$��v�n�,>V������Vx��'�������
��~҆��)h1�'�d�w�1�Uq?
���\Q�n&�<''���2D���=K^R�<��Ot�޿�!+���k��o)����4lF9����b��@�i��H�r��T�?���\�騊�e�8NN�TI��E���������Q�x���S�~�j̑Qg�!��k�~�u�^��~��\ �;�5t)����*u��=�%�5�?!�|��z���q���dvQ�[5�撶�Q�K�E��s%S��j��dV������]�3�߱ݳ0����u+H���-I�.��h�V�"۝��&NP����DW�'���O�D���/`)����Ǡ��n'}���<�M�<8��	����?�8J��n����vD�!��� �@jlF��F�T-^-��a�T�bF0�5��x��ӿ*��~\�o��M}��|��L$6K������;��	�e�g����w��K(9Q�z� =�E��y ��`;�����a:r���&T���En���^�����)�k�P��%�
v-(}B�'F}�G~ȟ<& �j�_j��&.�R�M�2d*G�����Ɛ�6��?}��;���>�b�_ �(3�h��^�S�8�S?>���&_���/5�W�
}�sZ�8�9��/��s)��_��_���#h�HN6�PȔ��|n2P�q���&T��`��s���NOM�U��q��٫��e�.���>X��X%�&"�^�MB�� �{6��L���%�f�\���c�ŵNOB���^B�	�����{iQ����<�l��P��_�0��T���g8�O>��T3�R��a)��}�K#�m����+��#z�����4'3	�]�-��_�t-�{����M�E,��+��e`w��un������PI��������Y��u��?�n7�U��Km����?���~�-B����<���;�~�~����R�d��q��矣R��D>�$��ŐI��FȄ�I���p��}���~y�R�tt:�t�߄5������`�	ȟ訁2�wc��+�u���$�����I����������\����c;��\ur�mi����K�+����o7�w���,���c����0��^I!��n�M�����X�O8����	~�ء��.��PH��G� _���).-qLى�5ùLo�+��Q�%c#'�#ΰ��U7�Lw��s�I�L�Lղ�����7��aǯ~��r?Q�gS�5i|?�� �}y���z_��^=��F�p�)T�6��}tz+�K�)��g/@p��i�qB���8>��	P��:���	O.��ZT����2r�5���|����+�|��_��n��4h[�u�X�ϳ�n�폙�K��t�ݒ1�꾹�[2�tM��F�� $�)�jܯI�kR��Eg|Z��B#�3�o��7q#~z�}x�w.�9�ib����>�9��I��.�b����ۖ�Kx�O�RS]��Ķ}�`d�~��yV$��IP9�r��E�{/c��p��B	��Fdo% É���P�͇��y�bɄ�=2�`U*l��3���M&y��������j����NB�.g�f���ӛ٫ObH&%ނ������j�w��ÙͽD�>O^x� #Uև�5�d��V�71u��cK�����}�Xh��x���j��{�cp'u5��k��I1��ӛTG=��;�U�!��l�l���h�{s^P�L�Z��x�Ң~��I2�� �<�L��K�k�
��j�_"�!L�����-�D��	/��Ke�>gq
�l����!�l��#��g7�:�ҾT�zs�
c�u���Hmpa�4���d��o�yo���z�i���3x���?A@�x~9u�5�3�A�&�-�H'���v��8z���u�q��_e�?,c�>���R:+"���_&!��1+�bV�4�Ժl84>�l�x�~u���.+�/M����
�u�",�R��7���\���ׇk���oN�� o��p�ƠJ(M�䦠�_ek��]�bZ�#�j�Iˣ�̧���RG����q�4�7,T��ͭ-r�~\7`Pi��%8U���;�������P��Їn�#�r��<����؃kK���N����3�,�1cz�O�s^�y��4s�%[ՍKN̯�i�rHf�R��.�����jjj*�8����Y؏O���Q?�add�j������Z�U��B�~b);S�je��٘,-��Y�b����Ӯ�f-cۃ����đ������;�]�AUN��ܼ<k��b]A;��KnW��uE�n��O��o�����L=�%�94����uxտz,����O�X���c�$ hk�W}Z��[V���8�᳷���ݞˣl�o/~���_�o:s�1B��mD�Lƹ>�-����O"�Q貲��[�T����$�;����L�Y�E���l(�5pb���E�Q��@>u���-�Q�m_iAwz����̊t��Xc��	+��%�MF^��X��f���$�4�,� � ���(yR@e?/M�����c\�w?���ɢ333&�.\���.�n�@��8�([9�W�#��#�í+N��J/����'-��M�;����SC�4��a��N n./c�끦<���ۨV$��p�ȝ6���'�~��_>����{�p'��	�&C���5�������������	Q"T�0���궕�[%/�|Ge�N��P���k���t�����-���f��ne^�N{��8���r�T�T�z�h`p�zo�X�e[�͊!Fո���g��)�pR�sXC��R��SW�j�n��K������g���L���{n�6����}�qp��*E����/�El3��ҰgO�q�5��*�w��@Q6��wv��66-�����M���k� :�G��[_i*�P6�bx)y��<���\?˻���
��)	�`���j�d=Y����Ƣ�GtI�n�4�#ܝ7J%�jp��	a����w����g����:��XJ�T�ݜ!v{�B�q~<Fqo� :�+诋��9Τe^=����h ��^�'}y�%s�A�ӊ�l�����+������s������@<�b�K��L��Z�$����D�/=(F�{�e[d��PZ潅]2ɴ���477W޶|G "��݁\!8*)9���" �4�@`3�Ck�;����sK�<PDdޛ�ٛ��B�}"Yw��T�4Ҍ��3qI���d ڨxߦ���Y�#̀�xWPP�����&�_��y�Һ��A��#�x�SL��轝�Όr=�7�i��>��Oܙ�~��hi�q���DX���`�����C��·ӈ�zr�9�+�|�x6�4��]|ZN��A��5 #��/o�]��3D���_\�4`��9�G�8�h���厝c����l�!�?''%~��=4��6�n"�dм���r�-ߕ��)|-y��W�_!X5�� G���h�z/V�ge|b��;��GA�9��V�4���oye��W���c�X#�y-�tg�$v���i�ţ���o"/7��뺁�����L-�s��k�ѣr��Hn>U/p�C6xy3����mBh t�{�o)���Қ������]��5)�V(Z1���ty7�"E�fC���p33g2�O�0ۄH���8Z��B��/�(nX*zM�~Sj�۽��H�.je����oO:ל�_r0%���u,C�1u3{1\�⏌��h{����NН���L;�G�FV* wθ��I����$��;D�Us�^-�-����/�c�7'#EeX�8��:{��9�{HH�h��I�P�bS�+!!���@�x����}ܫ|SN���FA[Ӣ[!��!ؠ��� �7-�{k�X�y����� 	?a �r�"�:݇�}��K��T����RӗJ�c��H��}cz��k����}��M�b�x���E�j�3���Vf�c �|L����ݗn[K�*gW��Oȝ[#W����R|q�Rз���q+4��}�Ri���M�6ŽU�`X!���d��D+�mM'R򔁷&��	����5���o``�D����O��+����U��Upے$��h*�5�>���p"���Y�As�N�4,�n�'��;����:ޑ~$zj���kZ�1#7#K6kA��P~ Nܿ��W�UJ�"4,��Z_��꛱�_5l��7�nN}4����$��J��q@9q+�������͛d�?�Լ8�(��"��`��|����ؼ��a
e�2S�^̧�������$n���\�B���P��X�jӕ2>ՄP�uE�Υ�o��%S&z�D�qqj"[�����;�؝NӠ�HӝDI�B�h��*U��O����D�h���*���^�܀d�Vcގ:?kmU9M�a��Wy&�|���###��u�E�nI�X�4wvi��M	Zv(��,\R�`0�!Be4T���8�������lzF���%��e���s	�	Sp�%/L��-�`E�~FӾ<��� �����0c )ZH7��M�6<nɈ�rb(�id�Y�"r�/cOʷ���O*�8��醌ע~������ﱦoRR�w��c�z���B7�R8��1o�L� �w�;a��s�؇�Ur5���ߺEl%5��"����=b��V*`FJa�-sc�b-�&�����5����&>�x=_BW��C}�<���\��HB�Fp�_�D}�=I��/��Z~�:}'bё���|�wR]	�B��� ��mZ�,%�����a�Ґ'��D*�m���OE�V�'q˸���T����\�����&��QM�����кIic�rJ���M�yyn��*'�U�\_��X%�eߊi�}��m�?����[�t@8���~o3�@QG��h.��_6��7���oRӤh�����9��8Y�aո� _�A7�ͽ^1$��p<�O�W���ƌT�����څ��&͠�W�������mT7�Kn)2�4�l�ecOx�@  ��s�vm0�����I�Ҿk��o:H��5�����6��q�@�#ťi��4`Z��n����C�%EF������G�l�l']}��d���/�U}<�����cw��������U{\M�׿�~Y_�x2,�_𔋡�K񟝝VR��ԗ4m�{Ct�7 K#��uH�n�w�`4�l�]u��M�ai�޹:M/;���r��R�����D�S�:!kW@��_ɡZ^;�|��hP,&+{��	:��/��	]����ckhc�Qѽ�݁�F�.�b6�x��
q��ЯL�v1v{W�a���#���{���G �b�PV�B��]�"��A�|Ⱥ B񺾾>��⮇m��9HA@/�xi��:�L�S���ٞ/B.gl�\��[y��	�|�i�Or��7����	$ot꺝T���jd-�=��K�K��_�� 4������K�����8�h��cb������V ��"�zc��E?� �#��v�ǞͨY�UC�������W��3�/'���7T4�yx��S%���ϧ|��<�OY�'XM��J��4�,h�Eq�,ft��f��r��=E�9��82��Tb譧��M�EfT��y�z��Еc�Oݬ=v��6�rB�6�RCzZ�]k0����^��O����g�2����6`y�]��{N}��d�����I�e���76�&9��8M\<_Y��e�ș�G��70�*7��r�Y���^����;B�@2E�L�֥�G_8�)�!�u�� ����"��ȋ�ȳ�704d�le}q�p��}5��*��:��#-�U��dH���/׶x5#�m�j��ePvp�~�^������ʞ�?_�mT���FD_�Y q�=����.pv�νRǡ�k*���qh�@��7�)'� �N �ܪc҄K�Wb<J�Rxq˵�T��\uJ��\o�=Ie{��t��U��;LL�C�KK�3���;���z{��r7~�1
V	������f�쬶��M/��C��A��Ȼ;{K�y�fu�,�(����\m��x����=��24���n�W��O��L����!���ì�����BŦ�MH�� ��aŌb��|A$X�c��AD�O�J��_�7����H6��ɣ\M����Ư���-w�g��	�J��������QqqqD�Eč3:���)" �/�KcD���ئݍBO���q��yHө�dp�����c�;�|��n�y�#'��*��<Dp�2�-2�KI����b���?�^,b� �
[ow�����Z��[g����R��Ȍ�����ʢNJ����^�j�\��[Zc`�L�_]��zY`ǘ�t�p����_g��_�z����'��r!�_�{
u�LdV��7�1&�����S�S
�������������ӯ~���y$�0A��Δt4�rl1mlQ7!��co�]ZZ�f�����Zހ�^� B
�l<ѽ̭�a�P���k?
�z��ʇރd��NN�;���mY�FCą(s��exc�����h~qQ[�ˤ[�Mn�T����g栕Uυ���o���ud�($�vk l����:�N��J@Qe��.]�|99=]W$����|���DS��Qc�hzr�D�]��hO6F��	O>�U���P&�l����8�"��⁰�0���m�,�|;���/�Z�hި,���&�ȴ���I�'@�p���>:�=�#�C? G�I7�c%aWc��)V奒v
�3ҤLI�s��}K����o�d�e��3pyW"�.�Ąy��Ӟ^^���N���8�uKM��y��������7>~��MćJ D���]���f��2�kRf!�^���� 7Mز�oda�o��P������31}Ɔc#"G��ƞ���T&9��Li�A��]l��1rk�s��j$�␬tp�2t��-�r�-e�yόx]������^F��2�PE���.��k������|ۧ����~��!{){<5N�b���^"��k��m���c��U�*�b���P���Q�-p��e�n)����K]R"��6z�7�~�k�h�`c���2���Ә���̫xh.�Ю�����%F���ݲA(1�e4���wǴĥKYfb�%%%��f� 8��(.�+�V\�~ְi5�E��-M�p���z��r7T�0����q�32�w�,,��A�>�k"�팩���'8=5E��K�SwvG�t�ŮG�.�Wpx1ܯ�lV����"UN�Cr�����;Z�)~�����Tn���f
�~:�pϦ��>�@�x�"���8��A�'��,s�������_��-^��-������ew�'�O��=J�el��/�a�(g�;��7]%����1޸Rw]��E���&2��E޵¶
	=�1X�R����������e�C��#x+G��k>3�$9m� {�����ON�T[������~�S�tjj*�O������/�>l�b���|)��^sQE��Ǹ �ݑ���vz��!�[:�bb8T��������[�I!����r<�WUIzz{��.d�(��I��c�^�1��ֳɟ
�<y��qc�Tp]���Znq���1z ���O�Aؑ%DО J"�nl�w2��DӄF��@��w-Y�!*������[90��{s\Z�͆��� C���*�;=/)�D������E�5P��=h��q q�ҋ�"���~t��!�D���M)�x /doo�V�@�.r< �Y�W���!^����5����e��_�Z�O��w������{��t�ݛ�v�-�!J��!1a�����ўW��A���� gY��J�Wm\_�}�8�����`uӕ�e��l��r��j��L��.h�Z��D��f��v��t�q�6�G�*��D���؆w�l���C��/�k�.�~hȤ��"=���O�&�iԛ6���x#>�����+T����y��D��ŷ��Y&�<А��^�l������^����U��cR��|Qi���0U��� ��wd!*�Ǿp .�����:Q�L ��M�g�oVZ.,�d
�P?%m5��K�3�y����0�qؙ�V�9r�3����0�JgQ_^^~�~�X����is��n:��N��R6�PP�g	�/��Y��MNN�]_�8K�+(B�E�h���7���x����*�2m�sxe�����!��$w��mn|�uϘ�M(�;�D,W'�� �@zY[��_�wN���@�9��z�Ys��EDp�))����Q �� �Lh.�]%��.�q�
�=SPÔj�C�����}��BPCׯzC����ʰ�:�S�P�� �M4�G	���W�a� 镍��|zS�6����%E/^���˻��LMyO7�m==tTF=�&��ާ{�ӂ���^F5|�c�����4Q�.���tQQ�d��a���π��|`��ge@���t5��O��ry�;p ^D�Z �����v��6@6��2ǡ�n�:�2H$ve���uPI0���
{�1ީ �Ey�;��񩈨����T!C�Y�+)u �j���X:O��1��0�}Y�H��V[�����n��E�ʟ�t�U6�4����
s'�o~yYW����8�xc���##==nD�)ej��Y� O����@u������[��;J���Y���s�������%�&o��ء~Wf��}c<ژV��ck;���`�(D/��잞{@��׹$5��N���-r�L~��D^��f^?�i�i�A��)\=��!�]��n��qv��w `���!�sXl����s���lK�Y�Ԉv(��
{�O� �oiъ�^z�Jx�[�#�|P3o���jD�S���bccc�蛪]�s5��!�����A�4���S�yvpyY����!�ur���|t���IA����<ѐ�m�����F�����B�J�?(%��H�ಗa>�)�*��}4bz%�F`���q��rt$�27��v/).^�tn��@n��~��n���NkG ���n��?T�5+^A6QW��x���g��y�ƀs�ZG�Z�w�� ���q#;B�s���4r���� �e6�[
x�����X��M�P!����;��ixZ��7/��)^�O�vk��z^�Y��������/ ���1�+�V~D������C��ɹ�S\����c��tG�����s��/H>`aq�X``೨��7�7��w-A�q��V������ ����%�j�4���d� ����ghNQ镴.����J��8Hu�aN�� -|��@o�]�%�!JJ�ƒ/d#6�q��/��wou�^�Tx�lS����=��R'����� ���s�	H��#LL�u�l�	�'Bx�,Z3��<��f��v����I$��A�S�	1Kߡ�%��@��k؇��E�1Л{���sb|�L��� �A�o*jk?���| �ťT�c�ةO�Ү/w�L�q(ѫ{�iy���nO %�OI�� 7Ź��c��!���&Y�L[@��*�;a�tl�N��A�ɞ#���r����)�V4'�<Z�p!B)����K�f���F{''b��\�
��-/��PP��(4P�m/i�)P�P.���Ǌ󤧹SҐ5��mT�:�b��\��~I[D��~8��,���,��F3PL�%���.EX%�coŋ���W:q��0E�T#���S
4{��/䵪׼=��9(���$A
I�UO!��J�i8xx|\,<��t�(@��b���C�"����&O���}��50$3J�,op����@���ֵ�Ѧ&�<��2ẉ�Z����t�13`t�W�Hũ�����Cddd
������\�)�|9�9����1h������^���� �9�PX�xɋ*����v��vU�p�36�ܰ`��nKHHȩ�[�	t�P��K� 7�!}6~��ThEI�n޼��cz�~pFt�V���nB�h����_���(Ͻ�<IR~��8(�|����f`�������i:D�wo���䲒sq%����\ƞ��sAc���i������\D|��{���8�K�ƞ���\;����Ob|?-����i���҇]o�x�>l=��az[�B��.���xs_?ߝ�}G�e�[��Q|��w�+���w@�ކ��)���	��0�\G9�'mK9��|����~�	p0
p1�䨼�z^=�*���ɐ��K�L�Jq'�o�\�)T:Z0�F�3������Ŗ}�X����-5��=e� HUw�`��͛)MMʴ|�(�?G�~UN���D+�I��aB�<iD�8G����2 *hOEI�400�O1��Ki�L���Z-R�S_�~G�5(T��rrr�W� ��w��%̨U�`���]�.���l��˴���g���jM��g��Ѧ�����_���R+`��K�y'n���O6��4�E�X�:��x��ld`Z�!!!��Â�G.+(ht��f9S�U�d:R��������yy�v(	u��:Ͼhn��՜k�+!�QP�,Z��O&�[�>⤣�$|}�o���m0�������b�i@�-��j|�e���T��0������$��/������g~;~o	Zq����c�}JqG_<���Հް�٘&0�V�8�bu�W��G�z������V��@|ow�߀J��uB����:)���?c&���mnn��I�(#�J��ٿ���ټ�ѧ��ӓ���pd��U��S:�3f3��C��n���L��MBB❶�|_\)�Х�h�(���6�����(yo�q�	N���h�.R�&B�t�͟��?6�;{�l2 <ކ�v�@����S��WF#����JE�m�V3	�4�x69�=1a��fϕ�kL풀񯮮�V[>L����Py�2�\��:���L��{��j���V��W��o1�T����~�t��yb=����,JS:�	���M��K
�G>���?Z�`5P�s��t���i��۩���?�x��B��%T�W[���g3-h��3ʚ(e�?���ld����#��ņW�^�sE7��D��'���G�����vZ^��I�1d�8	%�Rb�B�e����2~o9���`c�&�z�R�ġ��bZG� h�{�H���g�&#�ֱ2��i|@�pf�j˶���a��]�i>r%ee�Ui��&���-��^Z��2�-�~aZ�l�c*%ݵ6Y�XU5�.XڀKv(�� �,��@h���3E
i�t�����������?���@ ��(r�g�_k@���;9�,��ө�<f�=��03�i���􅬍|��5ȣx�y�6J����G[?m�|7�l��$p�LV�Ł�)�aXxNǱ�R�4�.3Te�Sq}Z���~���Zx�,�-8�^�~�P�gRISmIG#�+/S0B��hD�̶����9� �Z��m����G�ITە־[]j��Q���{�׮��v���ԕ�ѻ�$'4b�7
W�Ҽ��$gLU܏w��\�a'�ߏ"HHJ��8#^�[b4�V��-6���Q޻�ߌ����*ǡ�H�y�;U�e��o���q4�n������ݘt�"	�yT���C�S��\��}���l�}��{t���ͅm��i=Gtw8�y��=ȴ+�Rc>��J�����x���#�wrv9�s����gU14y �ѥ���Bj��oı���Jǵ���<��� ���9w�<i��D�
'Caaa��������v��r��.���T`�ƕ73�y��i	u���o������C#,Nk�k]xg&�_�p��y:����bQR�e,�R�#R#�91��4!?w�r�|Cãq5���9uuuh�W}�^����?�����Յ/H@��F���E���uA_Hw�bc�nς�f���gH���0��/�[%ԁ�D��TM׉�HA�=%�n��`���`>*)3����e�HN�����������
x*��2w(��Rc-?Z�h ���S�黾zU�0��11F(�7!�o��)�Nd��fޅ��
���w@��,/ȣ���&ct@�m>	9���"q��h�2��_�:�	v��+Wtz�.vv���f����<�H���RM��898���J\�}[��⌡�˷�a�u� ���V� �ҩS-bo}�� �u�.s�֌�+6e|N�`��ÄW��fbZ�Fa߽r&�������b�7t��������aȵL�Y�L>����ձg�}����v�4	p'���EP���"�&S2�zG3#h{��W[J��lii����r�����}K�jM��  ��@�p�w��)�W���7lQ��v(@�4�U&��� YlG�0�����G�/7����
>o�v�Ci|e��zp���� M�r�<�z����P�����u�@���HM��v�=zSp�F�=|Í������ �@�p�T�U�_v�#A�om��ҏh_lT{?���z.g??�p�׍tٕ�:P�9 ��T��nad�U>q�C��Y�i�C������^_��m��Hˣ~a��1�=�Ҧ�B&.�Smn����oRS���3ihi#��L�*�ܡ{��������u�7�N* ���^��D/�����������֣����`(P�1�}��[�&������?z`��|��*�0���пvܤ���z��:���.%���.<gn��&�Mw.���c���z�5S�}/Χ�Ӕ�PFg�br�-Z666K�KKW��8����ϟ��o� բ�c�;`Jt�8�m/��M�>����cT0:%=}PM�񝞉��h�ʓ B
��[:48�4�!�$3��\ -j�4\yu�ݫ~0^�&��նP� ��Ÿ���~6SŧY=,w2,Y��<�6 LT%;�Z�B�R���Xy�1�=��dO����S�e���S�B=_��t@� ��Sox�X+�1@���VQ>nNQ��7��JUϧ�g�o�M�,_L��
_<��i��'�
ڈ�8>>~U�|��X\���f�����&�t�y�/6��}�c��\^� r�����{i����� ZЌ䥤��I����^KŦ�&�R=���{Z�_&���&d��� ���)�<�Ī���:w �d�Ps�s@��B�j[��I��!�	ך�*�'�����Qr+q���E�������X�Ƨ
PҠ�9M��_`7m�����y�7��MZ����K-�4#^GRu���LY�ٛ�f9ݐ�*+���xwٻ��(xK���+�:��\g���%��WvP�3�x����E�G�l����[��3� �1�k6�nᒎ�2u�tW]�2CV��+�������K��>p8��2o�C�C�95��Q�r�i\[���,���0���i��� ��C��\�1�l�9���K��ɨq��#-ҋC�cz���}AW&�����կ��&_��S�d���Ҽ�&�o���ή����6���Vɹe���[�U�{|��5��ds��v��L�e�s& S�zՀ 5����p�Cbz���&&������!JJ �O����~�q&���b����G��`�xs��!�� ��t7Wz��B��`�m<���~�$4f?�-���ɸz�N�+��K���j%��s��_��ݾTt�z���' ��EZ�,,�&l�A} ���_ s	O�1t����KR::;��O544�������Y ������ɩ��[4M���J����?@L����`l��#LH�����Ƽ|i��Yq�Óϙ���Y��$�0�+����v"���ƆL�$+�\9�S���؝)J����� O�V���J5�Q��׼�O?�C���SDw����-���*,.V���8Ӫ�_;��k{9�����vQ��N^8��� R
�O�UW�+k�鳌���?rRҖ0�9���`"�FGU;J�M�t�GLR�#Wkԕ��l��������X�y/�.����%A���[
/�,��-���+2v�j*l=҉P���14��ɩ5���{X>(ܿ���KkF9� ����wr��
�r���ݏN�(9��tߙ�`��� �{/lXe;כæ��������>mCCL�)pQ#�!��
Ͷ���:�B�o}��W��r�c�F}���ק�]��_��wtp��4Y����t��ͪ��Z�U��UVV^�b?�D�Nk+?iF���&�x'�ȑNk��㘪+���  �@��:��O[�i?(%_����ǲ]_�r:�J�ȼ9M؊��=8*�!@3�s?����nY��|g�&�JLVU�Fj�(��L�n>�B��d�X�����c��ԑ-5���� ^���[[�,оx�$��&���i䱦�b��. �wYm*������ ^�z@>�M��1)l�f�쾂p�
z�����?�۸�B�E�4$7`&���j|G�k��L)����A�gg����;�w{�$����rr�&7//�6���س�4�o'�mf@&<8��H��CgI��0/B;�.�>�'w��q�>�cXc�|~���?�T	��n������'K��(W�ِ��g�On^͈�rn���C{�`~�=ei.�rZ�C3�@O��`Y�h�#���Bx~ء��K
��웞g���)��4h��T��*�@Z(d5�������������Nȕ"�^������ni��>����j� �\�o�(��i"��7>�z����-?ڵPOY�Ӥ���� R-)9��,��cm���]�����i�hj膢"����#%�fɂ@�m[w���уX-�]��K�n�v�iT�OaKspd��+?���l(D9���ч���{�
򝾐d�Ԡ�X��;%N���q=]�2���w>5zv�������O�
���1�'~c��靉��;5΄(��h��'�����{�)u��� IZ�t�ֳ/�*1z1����_���s�%�A�GW9a��]���"�����X��о��"%4���c����Ug
�d�F�X8��ٳl�l�? _�	\�'���¶T&����M2jj2��^�Ue��S��]m����y��wX,�*V8�`q��6\����\@��+�q�s����Yޢ��?]LH;����醫�]z80�w�E�Y����1/�?&���?���¼�ؼc�"~�oO�{��Ͱ'�SSS���z��
~�ѷ"�ۃ���ll�L�ʧX�'[#;�i���́m���2�tG�/�WSy"Z����I'LՒ��]��I2e��[KE�rV�p�0SQu��d���sl��1QQv�C�Ug����z�= À�&C��ؿ�HVm<8B�@��6p��ޅ<{���y a�� �����Su\Q�Y��C��\�J��s�&u[A<
^�m��2���5������V+_D���8p�OeQ11X�.�ح�l����L������)==�Ψ���{�@$X�l�5b_: 4�ᶓ *|�N���p'!�.��Mz�OB����k�x���DQ|��\�fI�R RZ~��Y��Z���Z�l�ߘ��-�!�D[ ��L<��Km����S3��w���Rƾ*�!.�����?���F��m#��d��H���"}��,� � ���c;����v�oSn����������X��'�(��A����]�o"��?��y��ΜZ����m{g�_���^���C� (ȸ�rF�OF�b�u�����w�����ӏ=6փ��l�8��!u�7���o��4�&Vt]]H{�6%���焉�e�����g�΅����3���^�H�W�H�uj��|�<dj�!R������s�L[c �Z�,�b�X�#�ZUŵ}��R.p1���'�m��u�3��w�uI���iۏ,�g�P7e���[��z;q�ٺ�C��(�1�pzH1*å�w3MHx�s��	D�`YWA�y���ӎ�d�$�����zw�bTt����P��4t=�dp��%�l�.�DaΨ��jﮩ~0���f
�!�BBR���H�[��o-�(�o%Aqy���m��+��O�w�H�������fL��zL���20>�o��|��/Y`��|�P��0�����Z��f��{?aj!��۷��AL:n�	��4a\͌ �l�����Ù�9_�_&�O4Tч��(��q!�P�������\0>{(�������d���9)(�88/���#��'�9�%BB;E�Hh�Ǵ�:�q_0��{���nw=Oq �4���a�	�(������wҟ?.�!~v�w�|���9�]��Ib|~��:T������U�(5���3r뒞b�v�HBE�ty�^h��e��v>%^p_~��}��T�TU���C��ͥ���TWY>UMy��&�.~� B��)-��w��_B��[}��w�J� SqE��YZC=�B�J�R���*�^�� �@�y~i�f``  ��'N�|��ܽ6Ut)��ʧ�=1A����:D�k��v�>�7�hO+LD��E�|6�cpg8;=?����x�>���?t9lK�O"��6��}z#{𶔂B	�l#����Kޞ�v��� K��Ъ �ot���r´��ў���-���/�3g�m�zz�FG3?��I����������.Kоw��-\������%4��yk��\9#�uf��MP���[+eu6;����d"����Yh?����
��Ҕ7o�o�Y�'�2�&P����b�ofr�����g�ܴ��M�K'�.%Yd��B������}&�98X��m(D��B�۽�w��ʉ#�K��h�9�cP��E��%��'���w�/����y��'0���\�%ȝ;z`��ʇOq�b9&�e8����&���Ie������u�T�ZX�]���~>P��߇�� �����4�Ml��t�srptǝS-t���
hzs;��UFSUԛq��#��obl��t��7\��A7�%��1�a���='_�sv7�53r��Fi�P8�B �c�9�uu!���Sw�Hus���m�m�3�X�$c�
~���[u$dg�����q��˹ߊ�z_����S�ůƕ��b�k����A��V���,:`Z� ��GO�C'��>��V����
��M �;TU]�����Ӎ9΋,��7�I�n9~|� ڠ�騫�qm�-�'�*�����e�?��*��uC�JC�@�Ll7��(�9
`����ō��~=��(4�F>����:��Z3��HeM�cX�D˥�=��ڎ�@����?���8ύ�y(�.�R�5
&7>��j����z@e)&9p����� `\aE�b�i˄L`�6�ٳ��
�����:Ҙ?\���v ���Et$8��Kg݌�~<��"����6kQ���c�Å�bWVW���Us��)++�t�F�R3�r�������Ri�d@�@�[���E���q�w�#�4�p�r�D����!G]p �ju������c�ys~�fV����/@q��eb�ImR��.�Z�I�Xx�����D�Ϲ�c�{	P1�W2Bg'�m����l`p0���CI� KBX��KDb����n\0�
����!���&>]�5w�ǘ�
�g^tc��7��K�˲�EJ��b*�S���3���iw^�y�ҸO��g�Bش�!��d�3�Zr<�%׿��#����#u�߾s�@,����O������#�`�-Y(��ɱ�� t�~�n�ف������ 3��rޣ����i:��ՏGʁ	6�R/Q�	AVz�E�qoO��G���bޝqZ�90Wy{x��LEmFo�1q���;`LI�C��0Ţ�E��J�P:n�Sȁ�zo��O�7�b�:z�9@4n��+��E�8�Ή���쒐�)�����W;��l�B{��$��=:�L��J��Ó��l*  n'"���<S\��d���.l�n�#QOh6�c:�@UR�	G��>��3@�	���94�2�A�yǽq�o�_���2c<}M}I��d���T���5�Ǖ$�	|��r��cWii+��:�t��+��b�l��R��'����s��\�t�j'����os��M쌕�"+��^G�gώ3e����=#�\��z�(�/~tEDR	i:�[�i�$��Ar$%��C@��F��a�����|��<�y��c0��'�^{���.�+�n6,��H�&<`���ef���%�g8���e���·���U��VVy��9��٫Y�ж�$$nBi߿k ]:��i>ٟz��I������ǒ����&���"���t�_���������B�;��6��iأy�q�(��/V��N��L���`���6��2�wq%�f[���b8PVM�ke�>��qf�(#ro֛���8-�av �=���{M����Z>������AL��r����b��$b����!�΢���[��P�^6�I��0H��Q����j�eG±�:�>3?�,��3�;����h����[���D��/]�Z��Um���O�j�':�f8����߮�lo��͗x�*A�F>�Cm�BW\��p{������ P�������k�NcK1R����@�kHX��~A�9����=��� ������2�n����C�͘gG��_�˫����(�P'^�h���T��m�C�
0�8���%�Z�B[A�!"�=�D���B�x"@P�q̖����J:ٺx츂��B����X#tycV^&F�䠬֍�!�S�;��GYYY��� �ҷ�2����*'-���2I����>:4c+`�L�	AvN���i7��_�k֧�9u?�_������l��Y��W�vy��8��QOOOB�e����0�ttt��ɗ<8�o�LLȞ��
X�1Ǫ���8<~��ߥ���'t�b�z����z��� �}P����u�24��2�!� `�v�̽�<wRQ9v�7\Qp7��?Q	���R�Ӝ��'�!))�5U|��Ho��4��@cr��:�-c|
t�ҐG$]ݟ�H.�?)ᷮp�;!S���=*nmƅ�}]i�x����Ŕ��w+����%��n:P��G�ˍM��c߾E��F��Ӫ�d���r�ZҺ�Z�Z����	�U�����C�ŁT�@�%XH�/ޮ��;�M�r���y���
aT�:}�W�а�"��ma�I�2?\]�,,, !BA�P���Ȁ�	P�@�IH&�A��n"ns���F�A�I�x�ӵ1(p�9��i���W�uq�OWm��9V��!��Rjv���r��)@U�x�,@(���\�mp�8�����@����oܳ�?<�fq�@ �K�2v��'�N+��^�\Q��*oK&�Vne��ayeY\�����go���|^ʈ��y��N�-�d��Y�\诲�[��.���M��?����и�q$�v��#?I�db��c(;zF/%�gWQA�z
���L���{g�ūW����ݞ�k[[�Rd���9��ʫ�)V��~Z����;:3�������Ά�����O4�����n�"�+�m����u2���W�*�m�O�	������L4���;�[��|f�-4��p�2�صc�j�ʪ��wPG�,�ƀ�4	�C���} o�Y���^r�����L_Fu�{����.=O_?c�U���n���K{Ճv��Z��X�4�_R���U���d%�wQ��_?���s�D�QZ�3.�"��No��OΜ�<��|21S�L��Z�_/�ܝP6��XH�`ך*F�����i^�
B�A�,=�����7>&�vZ�V��*�^��h�PL�-�bmN�M���?���DEE���{�c���T���[�e]�IQ�J�zx@�1gxX�1��[�,�OAR��uA�+�,�h0�L��h�S�Q��<�Qr*�W�F�w8��<#�R?�8]�zR!�����[�)�� ��[s���v���8��qQ���O��N��#�i�ݻ��Je�����߽3�@�JP8W�!�[��M8N/:<<LP) ������L���&x���^=��^���M�̿��$"2Yu��Ą�Y��?��}z�Ҁ�l���������zӝ1��UW�H�z0���$���l���/�=Ugo��Q����ý��|֗'҂�יVq�Eݟ�3�-6���PG����1�~��Ղ$����w���mRv2���]!��)ᇐ�P��*
�!"R�ק|�uNbb������b 	��V��t�v��=�qLW����Cer�jQ��			QO�
8))�T�i�5��ڕԶ[`U��9)e���mL�@/,|8��C�n;B�B�QN��2],��Y莁�09�)AMGW`���f'��i�,{{�	�F���ޜ�Z$Hm���z;�b������J�=!�p����DHd�'�j���Ƶ�H��.�{��Z@�c�'r�ʁk�Z��: V��҂כn]t��;v�p����}��iɣ�N=r�O��_/@����S��'W1-���E	��C�e�9�dw���cE�ڀ#ϓ��ӲʃW��������d=���J���|�攼&�^�M߬A��Ȉ־�
1�B�UTp= �2Q�Se���ٍ�:�G&��+C��:*�?l`��V�Nqsuz�Ҳ�����D�o��ma\E���*��8Pr�e�	���ee�E��MMM_����A��<��QE������zӋ� �!~ʗ�[��!��RP-@�
�]�"�ݩ��V��).�����}���
$Su��;+5���y�pO�S�W/�tcj���Q%����nEe�ʏ���r'���ԣ���>��S�^o�^!��o<?s�y��f�>��?�O�PQF�L��������I�Pхnո.��}���B����F	�>Y��	��' o|߷��}{�!��٢���3n��������.;Ŝ�OԜ>/��h��Ԕ��߳�O3����y�ECb'�,��6��K����a`����ʶ5�4�nX2�su���O�\�����즋�/��9���־�l��_��݀��f���v���3#{t�ՍK��	�t�̇ք�_3�RT�'@:�F8�e�Yߖ)l�XR����V�vHVx�zS���O{�0�o� ��L�U��,hSB!z���qe��I*���:}�Y�����D����3�!�\�w��^:w���y��!�oʕ����><�Ndqe���T����Y�ʐx'�<lg�Y8�y{YӺ�~�rm��LW�Z���[�c;}D�K]2w@���"�ݫ��qA�y~�	�"ɖ5X?����B���7#�˫[�c��}�:�ThKw"yV|��&lޝ����痛P˗Zy�j�\��X��/�S?Zr[�m����8Pkk���B��T�^���ꂧ�v�~��EI&�o܍�N��K��6�
M�<T/l�������b������r��I�z2}���߽�����J-�X���ez��@��j�" �
eîk��uEÇQ�II��֯G��ĉ5�8&
�ٜ�D�o_=��s��2rSް��bu[���@�O�e(h&ȜӒ�5���Vh_D���<�=�΁U##G�ʊ�%I�����	=�b�o�7|��[��J��¹;�}��Fq�5X;���O�Uu�}>g���|��ŭS`T�`ޑ��y45�cJ�-`�C	ؓ�$��:�"���^@M�z�� )?�Ѣ7���P�-5%�����~�_�� U�y���_z��ﵜ.�PeHeJ�����A�iO^x�e��'�����]8ɶI%�,+������p,�:a�H�>nJ�zF*CC[�����k��c^h����j�'�l�f[s���u,���:�&�P�5C6w�O&�z}[x�[��?78�\����}"sOU�:�)_�8k��#�`�>�u��3ޢ��V�̃;��y{��{Uhܸ�a�a�9�I��q"\���<WP��0��w����U�U)E�S��Ӂ�����ޥ�-:X6��8��CH�c{�N?�,��:��YTG
tb}F�7d���I�Dc�9l�0�F���yx���."�;6ړ矿�j,1H���������m�H�H
m@H�i@�B��ʚp��.iC�(�,I���M/���qGVx�KdZ����W�����9@���]���+f)���U�,���DB�\�!o�Q��{�wa����t�E�"�-�<$i��1�+Tq:��]hKJURc綜V��ֈԚ�&7�G������Kx��mI'�~/	N�F+Ey��䒙���2��m��j|�����W1��
Ub�bQ4���s-Yw/��k�, Iae�r
tG�Ǝ:�I�@�h�ԛ�~�x�Y�j} 8���2��WTĕ����w�6�H��W�
�����i���['�yA�,��D��ϖFK��j~�&���Qﾫ�_�7666��׳:Yk�Gf�H��/��w�s��I���	�z/%�50�+�b����{MNy��"A��6  C���QH�i+z��a�.�b=A�Y]�Y^su@h.���BW���P=�c�Q	�N\:�Z!Fb��:v�
�1E9a~�\5�y%8����9�G7h�g�?�jb�^P�d�����Hu��5��Eِ���_�v���$�.��"Zh���gUKt��xF�j���-<+/-u?�m��^��{h�j�Ĕ��kӚ�&Z&[SB�wvv��{�����i#�5����]hߘ�>�G)��܉pz�iQ���*��%������'�
x��Ej���B�g}0tM{�ص���Z��D�]}���">h4�^YY�qq�y��L��ǣ>�89�v//����P������j�o�22
���� � HH\JB����d�����i5S4��(!���sr�*5X���7.#���/j�q�YNA�]���U�v��E�[5EyK�����)�1U74��bd��D|ŵ1���]���iճr�UPئY�[\0Xj(����%��b4m�mS���_�mm�V����YD�e��&�U�H^�- q�����yq9���J���?`�]N2e��=��u�hҼ�JA���]P����M��;>4��:� �<�M�.~rr�����4j�Zu&�ۤQ���{��h�NG�t0t �:��ODc�dC��6Q@���]/�z�����-�8�������nW���g���YKC8˘�އ��dw��� ��sN���I�g%Z5D:K䑉QF�$�e/�Ñ���W.����OA��VTac���K���g,?��9�n�^�W&�(X��KYt?��Am/�}Q11B'<�1��]p���~�T�m�t��k���$H2�^��D0�r��}��~}{��&laڤ��f�*���������Pn�xb����V�^��\[ul��qQw�����Z���뾻�"n=����Ľ?`���I���j�]er��^�Cs�eR�T�0��h����]Y�6� , ���'Y��yB�.�@���
�u��o�3���؇4�,��L���wQ=;��S2�;*�!ɭ�D�NQ�?9���(�ڪST�(��g�#õ�v�:5z{�>�t5#W�[��f}X
P�@��Bqk[[Nks ֫���q����`��1����,Ho߿�0�Dv��[�@1��b��Iܨ4�6��t���&/�\���z���K^���٩�<
��8oV�x���R��]��u�W�b[3�]aQ6��1���M{�XI	�}Ļ6�� ;����\�.&�Gj���<���@Dt\eeL�Ie��p���8-����V��A�H�,�Ȱ������=��>v�(9TRR��יn����A>�y�u����W�V
� ������6o�ԅ4Xr�٬$tb���y��Z0��t��i�����������زM��,���.�/��6�D���������|��Ne�2����B����*p%�ׄ����8O*svͦ�/HKl)�5w V���Bނ���uuM[��޽�P��+(�+�&��C[�����֞�t�Φ�����
,�E�ք�L�R>j�Z?�?>����:�������K�Z�P��J1جƅ́���m���M��3H�q����I�?���8WP�h�����C*�clzxɘ*��1��u���� ��XVV�7o���5��)�1��/��?K�x4ϖ���<��V����9� �~�Z���mv���|g4}���~"���u?_ߗ�^��K2< �J�T���d⿂6�그�^�
�!�i��

Ớ���ͭB� m!h��~}�.�u"��yt��%�B�Nx\����&@M�O.]�cf�l��	!(h�� !%�k�C�$�XAɺ�y�9'Y�TM�_.�5�7iHf���f=-a�Z_޽?׌�\���W�kH!.TF�F�1�F�j�(:p�m��xuZ���q������
�����2��%���I�WP� \�v|�C�M����3.���		9���|%V��)�*B@@^h��M�m~^�G�<�Y������[,��C0�+@n"��MY�$�Ϭ��G�9�����s�L�F=_uޥu/.yP��-�����z>:��!$z]�ׅj�^ > K�%�>�F��
��S�|��kɃ��M���ad��K/1�:�âDu�n�on�0F{���F��&%K�^i��a�J�Ir� ,����l�S���(Z�|z�IiO���$�F[��p-*Y^~P��m7{~^���f)��X�����oNr���Ub�N�YJ�V���l(�����]8$3Į�� � bݽ��f���񡦥�7�RLQ멱h��{�
�.�qP���l[�ˀ���_�Hޏ����{,0�X6(G=�Ŵ���l�ymLTcv�6��,��˙���y�`�º��u ��Y��S��iZN..�Z:Z`�D3
+**^�[^y)�?a�Z9�	��������`%��$�6}	�)��h�M92-����^��ʴ��4�d_%f�>�Ara�е�#w~�F�	��B�
��v1;l��rH���1�s�^0��D��+�-��F��8�J��h�ài�~�����.��#��ad�~�Q6��O��:��4�Ǥ�k�]� ��>�;S�֓#Vih��9t t��A3�vl�ׅܥ$xx~���9��(ǝ��O�M��I����IfUn�R�� �Ϊ���(r�#��H��v����d{PP�2���M�}��0�~�@c���,9���R�;��	�}"�!��2mS�|���_�'�&�sn��^g0�Q�i���h���e�}*tA��N�u�`ܟ�^Z��7c�S��va/W��T	Ph ��,��v�0ښ	��F)��eb�J�~|_/�e5�.v�{Jd�u:Ql<�"��i�RZ:t��Aɣ�%��\�02�B%�BJllp|:��@=���67�V(���k=\+�&��r�a���$�k���#�G7N� �#%%rZ@�٫1/I>>W��G�ߛ)�\���6X,�ڙ��g��,Y�EMC�����%���.���c�KK�o�}�z�y	���	���a!���T�B^����M��D�m�eNj*�0N��c*q�k�	Mxy�U&�^]����@�T�se��K(�1���1�x���T�7h=1Ԕ��=�Y*��+&[;������v��%" ��h��l I�F=�C`t���D!�]�!�����}������K/��L��b��� � �eJ����ވ�@u��w���-~����l)��&a`�6��i$�ͻ����,ߗ��r��RA�I.Ԙb��eZ���Gm�4�L���
z�0�� -�j� �
wQ�ʶÇ�W���#�[�݉���Z���4��7�qֶ�����8�\�b]m���i����@%eݝ��(�UF��A5fm����Oݍ�ٽu���-�l.�hj+-���\a���ѫ��}(^Zj�'������A�b��?	u�)�s�d����6Pe��g����Iq�"¯_�m��<=� ����:����x���CΈ��V�����(�m�P���&F���*4U ��Ҿ��TUUE��v�hd��CݍXU���
�f�I�8�����M���4ť*���Y�܄\��B:Y@���G�� ?s���L�?�X��RHhi�@ĕ���TyF\�/��Z�I� �Qf���7���47��t77#��~΁�>�~b���D�������Ww��"��!��ʉ���Nʾ~%�*n�{>�0;��C� ����YZaA.����8��E~=/�����GFF�Jzaf,�h[�נ݆W�MG@'�+�R6޺i��Ky�6v%ͩG"5���_��!��z�l�ڽ'���a��q34s��o�������qT�P���TFM�����M7V����W��׼,-uǎ<h�ݳ�=�(P�Z����eB���$\�7`m)K��tO-��`�Od��X��$
�] :�W�-n��c�c��ݫ�,RS0��F(B�qtl�GN�.Du��LB^S)q��`.+%3)���c�hT��P������ge�|��J��L RԚ�EKlS��3tSSSs����U�5.AA�C9���0;>��bԥ.�E��!�S3T�%2z�D��;=��<Ř������܏v��3��H}\x3"֤��m�n�n����7�J�_]�����0��d��c�s2������,�F�PK�8���2)����?���Y�3�萳t�L�f�"Ham1�P��7,�ۥ6ܺQ7���9mR�����bS�a�����-�ȟ�#���Hº���N�WOrKQ��w�: �j�ųȯ�{��<��Mש����״&.�5z�l��K�׏���Q�H��G)��)��f�d&_����\]�[�t�X+���R��Ȓ��2�_Q���PC�ǚ�F����{;nz��G�J�Ê���u�_�4AU*1iyq�a�@��Ta�`����`r�sx���A��R[���T��tvz��x�%Њ��v���9��!"�F���8���>��&���}���h÷n��iO��P<����A�����@"��!ƴ��>;QȒ;�%�/���;g{�ݸH�!Rw�>J�N�<�FPsN���*|�H������(�L�M���	υS��.� 9�,ҽ%5��ͥ�i���)(0�YE���ݻ����]�Nk�*�L������FW����Pd��b�-V	��bsxD�0�~N#�)e��i/�jI���P��^I!#;����8wsn�fgg3}��_A9��N-��S�l��u������	P� į���������4�  �PK�&��jU]M-y��.���ܨ�T��]��3w��ͱ�&eCcJ^��������^A�Iu�al���!���� S�N��s �Rr�'9���hպ�u�v�r�n���Oܴ��[��¸ğ�@	�<��q&�҃��e)�k����(t���y_�]W�t^���{�n�r��U-.斜��6ض�z�d<N����e+�."]]�U��Ҁ��ZyEP���Fxz1ꨋ�9C��5'/A:�`�gr$��^m;�k���Rlw����*d�ЦA3�u^?�ym�o6L+��:�*���;�6�clq�֯_<�I$~d
�C5k�.1���$ �5\"��X���Jz�	�JJz���'A����:G/	;Uy�<h��Xp*����x���z]�sYu���]r����	�,Dq�^6�9���0���u�4�w��*X_>O9�&|L$/� ���Qh]r��bm���\E���|0v)_[[{t�/~�v������w��������K�*�DgM��M[�Dt������Xþ��Љ��3�7FM�SS����ᦏ���\}ɫ�D�sۛ����4ৈ�s^��6jp&����o�5�4���)u��X]2H���(��0�����i�����w|)j�.�@ˣ�z^V�Z@�[�s٩"o��<�_/ ���3���wJ�}��{���p����[NT	�c�
�g� �>�֟�����޷�dR�!9��غ�9\.��1��)|,I)���c ߁���h�I�`�|��<����n�,"Wi���}�q�Ag�X�0&��O����RG)���졹������ɶj�5�����әp+�_V�@B�m�&I��'a.T�ot���'�������(^ �k>|x�5��ȯ_��΀��Z�6�����*��T�%;?*wu;?6�5X����+�公*�.�w/�NMM������PGQ:���K)�n�w�o��D��@�<Z]��8GÅn�4����{���u^�@<�$k��xDLY��H�ˤ�W��76.HII)��D��)t�Lm+(00ӱq��z�Cc��#����▨{�)v��>�IQ�XG�O� �W w���za=]����l���� `B�,XNN�ፍ3�+�^[�mm����� 5���4��q]���V��;L�|(l)�Z�$C��=tyR�c虂��Uxn?~♜ @@ñ��]�&x�R��>Z�\�����Gu��WK��k��s�G��OM=���ݱH賴��}Ʋ$��y�w�T�1�K}_1:9p��2ь�R�G|��ܾ>��z��f9�G���,�׮]��#{2�!���+,\٬$�����bbzO�����f��ʄ���o�j��Z]��)]�c��y��*���[��5u�⫚���&2iJJJj���� jH)���)�Cx��t�A}J|�S�ĨB�5�*�&�.�,ӞR�i��M)-�<;�6Ԁ�p��� w�N�#�yR�a��v(�P�L��`/Lgڼ�����т�6�b=tNY��߫/��^�kx��;i���^C���.�����O�'|)��54����� Gq���X�0��T�� ^(,�F�w�:���[60>�����Z�#��L�Lt|~~>~�b��:t恺٩+q����oz:��	֝N�9{�U;�)@~cO�k"��5P(�@�tSp9W�	�E$tU̢��������R;Urguh���w��=.�� �~H�N���RF��*�L���V����=#����\1/�m`��	��{X��Z�'�M�3gM�bm7�*�+�x�F_w����{����J�����#�=M�Xr�s�R]�b���烙MY���Dt�p��E����c3N�
� h��I���-�^���&�ĩ��V�INd��-�Ւ�L���p�;!!����B<ِc\%+]�X�!T�F�d�����/]ʶ�G�N�>�Ú�*c&��#(Gs������ǧ�v--31l��L<ij��A&�Œpk��uВ����aR��5A5�2��ؐ��2l�!� �VX/�@VVV ����H,Ɉ7�w��_�y�e�4h'mnp:���KHT!��3��ط0ڢ E�sv���[gS�~�@���n��~t��*�=zM�����	"Ү�A�!�����E�ZZ���("
j�?��
|n�|u���&���U�c��+ Km�`�_5�����L�~(���+J�vo9��oY�O�4W�.IP��T�0�ң�d[|����P�V���`Ogܤ�aoб�J���4�. L�	��E���}UFB}�7�C,_R�yg�w�����anWyE���sss���RA���K� %���Kt44GF�'O6^��*:H
������7��\ �<�$�3�#�ohtTg ������T���`����d�;�7<�_p�k�*��Y���<��
'�u d�	�<�8�U���C�o��;8��nw`V��͌P`�B�{��7�P|P�ӵ�(W����m�>kR���<����]�&:�p�( ��Q2´�o޼%B�zy��!��H���湭"��ḏu��;��F�PSv~�66��z�Ӌ������(L���{��G'�Jq:u|½�Wo��mV�\)��O�����upp��z蜴UԵ�kdd���ll@(P\�k�R� a���p�}�JP�~��|P�k�fTL��mU�LV Y�,�&GӞ���c	<5C�i�g7��@'�|]Ԋ���J�"��h{e��h{��_��c-�3@pLR����~�_��5�"��B"�`}k�>�/m�r�W/BA�����u�X���2wƛ�2�7�B='�c��4�>��������f��������bu��D�䉛�k�"����RR�w������}ܔ��
nm������w���4�y�뷿�OH���}�
��(�0-�!^�Ͼ��,rt�qe  L���:��T�ϓt���Y�����W�s�	����O�-nu��YW��㗉�'�Uno�k��BS+�ٱ�������n�H�C�Mhr�s�)aD�$����	:{�y�T����ח����r��H����jWWW�C��^$/TI�]dR�V�0^���ݔA��.�C.�^��#�����(�����OO���R�Z7�Xv� 햟��j�FFP�Hʬ�tQx���������B�ί��<��0�#'��N�����R���A�<a��ˈ_� ����̌z�R��ޟ�����m����_��ʭ\ֺ�IK���[[rY��;�����w+�]h	��0�sm/�_$t�:IOCÞ�Ӗ��֐݃F�4`�D���9�xm'8'��t:�����u�R���,�ǉ0(?��ŏѵ&�#5���ם�����yM?ҫ4��?i��S��UUU�DDD$������qݾ|����S\X�S��E���	4hƜww轹	��N����˘4�s�=[y9晿.Z�UR���YI~C'��D���IY�����z�<�W{]�Q}���.3�'��#P��R��X���>��[pY���kh���&W[Z�q��?�Pow�}��f��H���u�89��ۘ'��c��Qr��С��sH�)��X@o;<S堼:>ɒ��x���N�#�O�X#%.�vrr�4}�[J�Iy&]SS#��Ύ4��p���]c;<rT������-&�ئ@��H��:�s੮9^c��)ո�,��к+A�MrvVN	��杒A���ec�r\��A��0Iӫ16�4�`���K|8]��o��X�5�V��RG)�=��	����4:1�oqu��G�� c"55��C��O�%�~�Ee�<4����J�����g�w�	JLk&~d���Dia��@�F:L�I<��6D{|�r+�N��+[̕�:��@A�y(��xz�ǵ��ǯ`0l�J:���ccV�sdR�<��|��#��of��_xh��&�1�Q>�k5!	�U\��〓P��N�v����-=����3�E�Q5�?k$X_�Ծ{�f�&�-P#�����ӎ;rT�z�� S��f��:Q���}��?�����y o'z����]bbbi�,
%�"qWB@@��t������q��ڵ?���]�����t�z�f^���o�7u~�#�![-pX�����>��0[Vb�鈨����|�6I^�g}ZF����^3�X�'%���%?���@;�Z&��%%�<�y"V��!���F -�-���'�#Y&���q�t5�=_֠��̌��k�tb�ٌF�r��K�p���8��Fbq�kpڲkc�KO2��n�����;��1WR^�b�s����s~~~�,4Q��6�k�@%�IB9�Gջ����e��:�΃ާ�&HO.���
ї��,�O�Qq}�Q�磞��n���k�o�v-�Wb�4���鎂���5c��Ҭf���Sw3 ڮ�9 �	�r8���+J�t����������?���51����<.��T�hc�25��w����rp*kR(� _��	�L�;R3�k�ɫ�u��g��22U߳���*)�L �����a+F��~Cߦ�\c�D�~�5CC�?j�!5'�>��@背�{�Ne������_�:�;����jIQQQJ۞!�^�1�`P����?yʡ�!��C���ˤ�66f(�������'���75�A���Rj���k��>ibk
���%�3SO�:���X�dni�	���K�=@�n4ʃ8���M��}ZM��t�}[)�Qک���:��"�V�S (��q&x�h����<�Ǳa�u�\������m��lQ ��}�!e�*�+�5U�$�Ӳeee�5d�IE��RW_J��1��F�`�y�_p؊U�o���T�o�I��S �-���� MM�>-�%��gQ&
^7  �6 N�Q�m�l���?���hdoFS��la����|m�&(����h�\$�'\!O~
��gąν_�<\kG�4�f˲ǣ8A�cc��~�G�\��֊YF���7�Ʉw4��΋���?���w+��r��;��=RXmI��ygP���n�PJ�uyttoM�/��[��Nw��z͸:<:.3�@�f'�� ,���\��?g��0݂�Knok� 0 ��(���D��(/�Bל""��G�0|o�S&�L��n H�x��6�]�]�D��K��O6��/	���d�bT���j�~���B�&�`dIP7�yID^������8��B"��)��|!�!�6�Z���E�����	?�y�ڹ����殮��3bOZ�x%�O'�܄�4dW����8��N�MMM&ו��2�,7�����׍��/�O�6�!�?{�U�Ӎ����13���������Q���D���PJ��:4jbi���N:�9��w�9��$Y5n$�{ʱ2�r @�4����g�zmx�[r���iA��y��fb+�
��)��[�Qr����c�o�j_Ix�ɐ�� ��t)���ߘ�� ���q�k���
X&b�V(�q<(xUQ��H+\�����\{Й�;+�󕦤����,���]��}�|иA~���
9���dJv��lbb�����j>5����d�mP����󌗉�|M%8�9[5U��������M�O�c��P������mh��  ����w��TѺ�������7�/���3Õdߩ)�X3��\K������+���S�h�g�H�������}v�=�:,���i�{Ӣ=��VewR����E�'�V����P��t��t�r�Ó�!��c�۝A�e����#S�- ���쉃z��kSR��īL��# &�a�&�I=����G��$�1YA�U��X�Z1	�R��y��JN��[���p�-�C�����Q
S濉w�D�٦�{.�C��o�q��P3Oyߴ�|����L�uF4����ޕdB�9:���b�8����"�%۵�����03{*?�vm�@�ę���2^s��D���p�LBs{�qZ�Գ��񍍍����[��|o�/�lw��M�5]_q���O�U�cjr]V�F_�x��2�SL���oZЛ9`�<$�BE�^�z�y��ʄ7�F�Z�'U�S\�*l���9�J��R�s��6ڒ0�����c�F"n=�"��;2����_��i$ҡl���k�-<���tAP����R���Iܽ
C?F"�9����A���snnn�?,b��%܀I��1N?@
���@z��E"d��ii���LPt��{��3V��>㓚�\��Y<��^�U q����.0�:���$��	���r�|�ݹZS8
�P�3c���_���Ȥc/{xxԮ��Uk��r����py6����U~�@2���]�ƌz�W:(,��TO6��sۻ�T�a��>�z�y< ULl���*�3��0\ɢ�����-��@"`�-�y`cRkp�1�Y�4la[ZeÜ�IhS���'_ښ�R�+t� h�S!n���#',f��߸�MGn��>Z�YY��k	�t(rd�q~]��A;\�=\�_��<�%��-`��KD��)s�Y}���8F������������;���?xˍ�O���j�C�R"����R߼�:�H���`��w�}�p�X��%�s�m~�h �h[U(aǳ���V�U8���L	?��$^��C�[�a�J�V�'*�~�͓��0b3��&Cr�m�ڐ=T#St?� v�^����#�0)YY�*D��ڀ=�?go7ra�Їԅ/p�����ek�ExH2hMڸ}���{�Y���R�d3o���OC�sG\>o8ס�Tt���6@)#
�j��"x:�pd�t�Y����V�L�J�!�O��}�Mf2m,��U�%:�II�8�7m��Њ
������[{{��=CjU�Ȃ��e>��t��j�y�{������_ԢG�5yZ��жR��IIA@dTR�7 &;�9�Y�1�� �¸�o炤��������)�s�M_)�B��M�p_#2rq$����ȗ�f�_%�b���#�����dq����s�!�B�_A���&���-_v���;J����s�
��r�?��6E��?nA�|xf��U$5+���$��Z����W�o�B	��[,<b��ҙ#F_u��"dX�F�Lu�&L�UiSE�-���хF���V�li����7r���_4���B� N�����z��A�����W��a8u�-4�3��30M{ذQ%�b�J��p�"H1?0��9��r\��k-x��	S�yo��=E�}��_X���Mq�A�ia�ez��%+�/a.%m�W���({���0�[ܤnf���w�I�W����I�����f  v6�e��o-�I�S�g����^H�HBw�j�?)v�l޼G����$DN��7�}�p��K囬����sk��u�H�"�| ��?�|���U�PD"�ޤxi�ono��$a���N��E�	������C7�Xqi�.��0���>A3��y���B��_MNR?�WV=���{�F}�N���9�~"�+@���<}Dw�iz����܇
�9���>ZT�ԓ�8`I�~�d�8ڨ?���I��MMq��#X6�R��K�3+<(W�I<�a���#��o�!a��X�Jbŗ��h�ݚ�3�֨��6j��TZ�ӡ`v��eE�_I��N(��"yA@��*�}��G�h��~��E���D4"
`��m�FN�C�Fׂb��ֶs��ε��ʞ�.J^`WN���9M�+�eC�j޽< տ]"�i�:->Z�r�끪�����d��vs���5"""1�u1��ML{����.��K�c9M�Щ�EG��Jы��P=65��z��AAo�ϥ�D.����w�R�q�# �C��]�����V«o`���;�(�8w�
~b��K6�$(�%.ҧ�n8�,r�y�F����b�)oVX]�e��wO9��J[_K�|�U�u����Y8;0/E�X0�I� '���X���������V�g;_�^"!����c����E��[�~~��֡�m��M㘦���tY�|z?9P,ֱ�tK�="2��K�0Ƞ���U=��1+�9^9�w)q����p!�����VhP���%�B�r�Ҡ���P�vT{ �P"/����o^���R�l�ɮ��:[������t�Ö�'(ׯuE([C��'�Sь±��*���Fq���X�ߝV�P����N���\I���MJ�G�݋MIs�q�L�Z�+Ѫ�Y���?��Ȅ�]D,"��M��[����Ƞ��� ����Ѷ���#��:�s������z�?V!�����FA�(l��u"]�z]���id�:��BC�\~/7�J|V-Њ�1+��p���������Ty����|��Ifb����4����X� � ����Ŝis����`Ͻ�-N�T�\V��l���~�lH��b�$5�����B�0~�L��+x���>��|�	hc����ٿ�0�����?L]w �o�?H�"e�
e���������u�Z$��"��ޛ�	�{�co�w?F������<�}_���>�纟�y�������B N ��0?�2A��:�A[j2I)E��c��!	y�䅬OJ�r݅�9+#eA����x�bI�[�ۇZE��V]\L�����!y��ȱ����/�0Cq�n��ϿZa��sS�V���i� ��(�����D�Z���T�I2H������J���ӊԩ�7�XZEj�O�N���%9�"�i(>�Y�>�&}w�Vc��c���ʫ����G��lm=qq)I=����F�J�X�?�7
�Zpl�U�����8?�U_�{W��'�D� ��.�h�4�A��[rW�v�"�<��R�55池��ۂ9��`z76uy������pb��Q�?������f=ͥ�t��Fp2U�E�������ra�ΠW5�z�����cV���W���"n��%I�A�G��-�N۾���%���|��g���ĒB���\���u�P��l.�Vc$=�
�3�� 2尨H��d�u���Vdi�w��9^�!����p�nYW��g�a�c�E��E����N�o�y���>6����aOq�Q�U���S�p�����R�K�&Z���K�N��rw��ݛ�6�/��ι�}@�r wKd�SU�����	�ˡs�{s�%���V����\����}��⢓0�mq�� �;��4bill�3*�%��/�];]d̹�z��_�6��;h���ϱF�����kV��:l��:�^b���1�'m��INX��3;>��}���'���N�f,(�P�������ߠ��|���oJ���k��e#N�.�����#�����>p�����F�)���:Ar���:�B7QL���g���)@%���N*~�����#f�����Z�&���Z�����S!EMi_���V:��#��Ag�*��l�*m�Qz:��Rݲ��?ǀ��Q�>��KE;��ay�S����_�����W��R��iR�}�?2�o,)��xa��Q~�������+z���,��	��U����f_<ߝ��J]��+X�.i���BEĤi��<�d�ykng�;�2��ZGV8A?ft���p/5��oo��ǲ�U'������s��q�n%�wwu�v�׌C�)��wZ�1��H��E1Sc˿L���"G�1,.,����mF�?�{Z\X0�X3��9\�p�W7a�Լ@/Ƕ��M'��.�|ys<��<F:�>sx�$���0��W��l�1��|Q��#���0�$m����u�X�ګ�)K���-���M�>�Yl��"�����m49{9�^�s��-�r�t��s���R�o_<ӊ��D���a�G����Z��>��S�����$��%a�����K�
4�Y ��~���hG���=� �Dٳ=�'����7n܉e�*-5�{c��I1���|����)ނw��5u�Eh�-/{u���� 3��{��9�H]/��Hmm����Oyo|0�ߤx/u|�rxq���UQX�h@c��������[m�:�_TI�>����l���H�s9V��0J��vN��J��3��O�U�Dd�]�u>��c� �Cq��b�{y�����+R@�8�oY�`&�٫� <��b ;�:�U���=�'�k�}��`ɱF�PS/2/�ݺ�<�����aX:���Q��vdU��z��p�CܡG�ŝ?sx��㎖��Mu�Ń�� ���(����z+7_����(��v5[[�����3��K�Ci���1�_XAO�R�������j�^�[��8�!i#h�*��A͒:[�����������\�e�ɷ�̈́�u��|�߽#�d=Y~��Q��q�m�퍌 :d�����&�ci��lb7�U��V�A���%l�$�-�����q����z|���:6��y�<�H�'C���m�l��=d�ª�D�c��KQ�����4r,m��	Y�@�t"+���h�2�����.�0:����~~8-�^�`�Q7�'z�_srڱ.>h�#X��"m�q�;ֲ~K�Z��t�,� �ǹ&2,�����\=�U����L���i����R�.����ݴs,�2��K�lw�˕ɽwܫK�71�&����n�O��$��	��)?�*�L4��HU�a@�P�Ő�8�u����?�}o���[���I4FA��
���z���d�uCܼ���H,�hr_#�����m��bF�o֓}i+7��st0�;��kk%&׳�C��х��J׊� #��S�{�[�=�RI:)����ʊ��5�FS�\�e����q縀�{`���>�Y��U��vS���){izs�,[��~����Um.o���~>;�T[���۷ɉ��w��ߗIWN,�����h��9�Gb���O�E]x翕�(݉H6K��'w�wF�k�����.E�|�0t޳?���>v:�'�f��?0j��o��7��f�z>�=ꖧ bk<09����AN�x|�&,���Nd����'�����<��K���-�4��)�	�W�g��'آ���쿲/�͞O����c���\J��9��B�Ky_1����H�����������:��@� �l�<Z���P�@��qA�`T��"���Ԍ�dVUv����P��Uzn�9�UzN��ÿ��\E�0�v9��D.�,
����Ӡֻx�w|ܠpHG<1]���8l�35s���x��������h2�O6e3�خW�p��'|�{��tll�k��B�w�7���[3�w:K�u,p��|������>TV&�;�����:w��j��Zwi�)�*x�X�\x~8L+E֐���MP
֜����ݫ�\=<�������?��A~���@o}}�F�G��(���D���
R�\���9�+֞p�+i�T!C��I�N�<U-]ɫxM�+������i	6y����Z�N���:��G���_�:¥W.�V����:Q{��1�@%w��%ӾC��o�|[x�0U�p��]�P#���l�bDDD[�ws��X�\*�*P���FFFzg��
�j�x�zOq�b/8|]������t�.�CK�b�VI<�&��0�G���<0_�T��έOn}�����B���V��3��EΔ/x�b����bxr����ҿ�<�ĒȮ������Ci��l�˰'w�B)�GG��]��������[�3w��wv�k�R��'�lj �yf�K��dp=�W
~n��ZhYCS�*E2�j��C��M7Й�M|]ǀ��WB\�7"J���}�)�]VJ�ӣo�xq@�G�d��`}�����N���I���iV`�ul�K�r�޶׺ �j�vi��o�ָ�o���2^|����[ZE��������3���Z���� ��0��r�"��LR�<�	�^u��ષpj�-Y���lfث�� �9��ڎ��`��>�ۮ��ԶuU��^�����$��:9�U�>t��ڏVn��%���Q^w��#��!.�(��z���	%�(f��ş�v�g6�P��x%T��v���kZX�}+�P��M�NP��M[b���'�(Ӿ%*�ϿJDd��ibec��]#���Tg8���n~�=�v\���x�{@�W����
��o A�3�(�_��g�ݫ�B���LbJd|�-��vt��距�<��xb]~|����e�����\���TogѦ3��Ȇ�x�Ig����dC��ً����姃�>�6��Jk2��� H�և?��9��.o��]C���"�鿭؄x��*�7\i�w^R��AG+�p>U!��̱������D�!���X^�P���._�?�2��V�-x�%2;��5}������ݓ��5���b�E+�E���hb�Ϛ^NKKВ���f\0}��6�g��2:��2)_ZMu�5�� �)�QG(A�ŧ�(k��P��H
���o)�*�Q'�����U?���������|�׆v����CX-�
<ݎ�^��3{S<:�R��ȳW]s�U�u�5U�^���=���ݜJ��3$q{ 7�*�,,�ο���&�7����<��Yu[��gG��2\��~�vU����Y��ӻ_ϳ����(������+%�G�[����e�fj�\�{i�+�E����{��wm�����~jjj3=��pq3�_E^����M�G�>ۢ` jW���U��Z�sasw� �u�lP��B���	�RW�;��΀����`�:	�����M�3�X)R��%�	$�Q}4�e�_�-�*ɫ��,f��w?���ԋ99�^�.���b�	`�Kߦ�B�Q?ֽOI�u�ڿT5s#|���}�{�O��G	`�v�: ���;y&ѶU�xcF����vwJj�]+t�� � l��v��hy���Q M�<j���*
q�]��F�Ѹ�,���=���WVV�:�˟���Dp�ͥZm�8P��5>ma����>3�A���#S�����^��h��D-��2�<0�C�^a��C�{�JF��`P��X�M�:)�&!�D��pM�q��_kk�Q̰˕�!K��˜��m�x|t@��'��(�$^�ځu��ۇ��Ź-1�����1U+�$�!�����6lP��g�l.�=vY��}�k2ds�=�حX�J�{��L�ׇ%>�
��>�BoSnpͶ���)1"���YT��<$J#�z��bуy��px�s�j`1Dm(U3.��rP�"��ݔ�nj#G�aI���e���/�c���z&C��C_҆
�-uL@ُ��\{K�~:|�C��-�X�N�S��˓�ޏm]V:�9l�=#OAI����+
���谪�����x��&�D\��ѭ,���V�a���C�Zk3 ���r���s�xǖ*XF%r&Dʎ��S��@r߇>�[���	<g|�]���r�A�QB�k&ѷ������WRM޽P�w��=��}w����>mGk#�k|�}��S:��؋u(�T���;���P�f	N
����orM]���Cx4وE�Wk�7l�1�yz��~��p5|i)�E�O\�CiX�OO������#�,#ܓm�U��I��A��,�? n�^+[Ά%�����,�����($1ٶqП ';{�z�(g4��,�Y���F���"mA�RHnF��񍍍2PB��+�xG-��㞈P�@�>L��P�:Q��I�7�_����W�,��s��ӍԶ>פ��'��<���iޑ��ɘr���lk�bֹ�f�9uy�kS�{���xMM_v{��ѝxt�kH�m�*�o�����p��?��2�lŐ��9���bKw�Wd�~Q�-r�x7{w[�n"�����\��vY��5{�Cȑ#�����~�_豰��1�h�@[�%����'�ƍ�^%���5T�Γ~��Y���E)�T�G��qJ����8�\)���'��d%<��dO�Z��ѡ�hh��������_���
?�8� �/M�&���23��*=ѻ|�~	�R	}~�άC�����{�6��p��s��U_��� ,�8��	 �,m�[XنN� C�xJ%�x�cϤC�xarR
8D��?��YZY4	���-�]�BYl-���k�$^<~:�M/�0�5�PDإ��e"t��s�Pz��S��&\��@���~�WYIC�̂�a�]eP3���?��{7�<Ѻ����). �>�#���+A65|ɜ�
L�[���7��Ɨ��3s�|�ʼ"Bl�X��:��Ӆ��,�A������������oҾ�UX15�H�"��uOO&���J󤨴�*3���و_U�Ề��� .����=�6�@-�Jш{�&��R��|ؔxД@ {�ǒg�#�9j3.���p;|IP���R�eS�+��p�4`���{�����0IC�V�N�D���H�>(�����iR*�9,��n����H8Ȓzp��n8��$��[�Y"�/^y?h��)�D����k$(7҇����$`�W=f�͎�k�x;���NΠ(t�3�Ƞ���;�8f�{3Q�������_�<��NW��zU1,w2C�f��������swM���~NX�?ܔ� �u���؎�\;Z]�f� Un9+;{L[�@P�"�P�m ��G�|ŗ�ķ��Fp2k�3]ݑ��-�ƂvqL�����n}6|�ݚ���~��IJ
��DӮMY��N��ϟF<7[��8 �j^m��:��n�ƌ�ݾ�bm�h&H�����W�b��d���1t5��
�u���._I�Y|4��A(vC"����ȥ.8�q|��[�HӐϾ26������Q��\��th�2^ޛ�>����W]{r�2�=u�Tv?'<��XJ4���`~�H`
�����<$�`�,�iJW�W���b��3*?D\ځ>{Se\1����� x��G �gq�'W}S8Kx�哙�4��&$q�����<��J���a@�cl �	0��8�������W zEQ��Hu*%x�fs����VJ8��r�9�;�S�,שO��7��o�#�4 �cO:{�^a!��r�KF�m1�?1�5y*|(0Z����9��n���.*��r�̠�A������:���qT	)�'�<����0K g+�s�p�|��3���`dPE����i�.���(١J�u�1	�:`jf�hQY�u %@�	�V�y��r���}� �m�B�abr�9���K���Wj�)�����*^b֢X���W�6U�,����
��"�=�T��m�!�<�KI� 5 ��98n]�)}T���d�W�2^�KxA�|ff��	d��X����bdz;��T�����k�~U��b83��F����V��)�]$#{"�QE�)�����h��'�\iDف�i�:@`�T]�u͇b�{�˰�������{{MLR�7#�A'���m`d$�,ыpw�EƵ�p��fO���o�%�&�� \�\E���s!��bO�3eX��0�*�p��s2A.|�|u����I�G+,�!:!��R���D�D�t���v�\ms��RG�Ē��б��`1��	�o�h��w��g��v�
?Nb���@~C�	>h�3��җ����K���v��=`%�F�@������/����NáYy���^`9:��WhC9�*W���~AL��'+\$ Ё�>Y�9=$��㸪7�e�JK��>\t�:�6�/��p�7!_������<����s@A�$
Wr ��Q]��)��I����u�.�����@�����s
�o���_Ck⁍�х����ʿĢ����vkpW�W����V�߈v�<[9���_/��U�K�5)�q%̊|�Q�{��R��ng�7 G�Ұ�ڟ`;����d|��ĹuH�umT�y�Eؙ";V~��(?�^p���[�����R<����%������'c��C��s�=�K��~K붠���&�TU��~�X)v2`>�T�Ar�6�Ü��>k�����Ү���]�ȓ1;L!W��yزǾtF�O���V$��5���	��Ȩ(J��J�1��Owܫ�={��:�\9������8�k�Ve��h�rG3s���N}������0�jm43�oT&�A��Bo���r�Z8���^۽=�U���G��߿}[*�.����8�ZR+��=�@5��x�z#� 	\����M���b����L٫H��oJ��Ûz������A_�J�R��0\��S9q���tzg1W�~��Suri�o!8�ψ	`2R�$.^��^3���XQ��Sݏ��69'�ݓvE�7f1��4�_ݪ1�xȯ���>pU�=IXa'Ш�z�0���5��`T� �^L���!ШDԫLp@nQKW���(����(��a]U�দV�v
�П�Ӏ�C�˟O��}��Jx@C/)T���Z�����Uw�Z��0��É�� �؃��[j�%�ԟ��l��&�¸ve[L�g�c�_�prq�c[�K&���989�B��j�@�����t	߅���}�~��1G�N@�g� �gz������[�h��!��x!VN|�m����ޔ�u��hPTgT=҄B>��Ʃ��8	AA�����&���w5�H2ivv�zH1���M���555U ���pm���9��W�������S1�	q�`��ga��l��,�uw��
8�@��d6dh�ki?[�h����f�9GM2g�SF#�^�r�}FF��Q���E�_\x454Ƣ	��A����Uq����,���H���쀸����I���,�z���Zw69nv���
�9DY�זA�3�ڟ���a|��X��Ӝ�@���?��S�Cz��|���4z�i�(<����WݍVe����p��Bn\:��m��p7�2L��Te��f.���5j��i�$�h�u�I�ߠ=�������9e�!ڼ���X
k�p"��쏬�W�I0ŨnL���hd�)�?����ax��юL����z��:nB����o<�l��Ms��j57�(�0ɒ^ʅG=f���R�]]]�S�p%P�*�W_��^c�h��<aUfUz���$�� ���<�W��|q��yN�eQPPD���:��YD�U@`��	� v)�8&�N�$E�h���~eZ#y�&�qos��{����2J�t�*}[�7���3O��,�]���g/�	e?彉��)G-Zǈn��
�Ņ���Wɬ��K ����qm�2Rͮk�����յ�r#�E�|1�!@{��@�U�$��ܱ�/�@Qr"�<���]+R��hx������
���Ӥ����4P�}N �4JNՎ���h����D���8q����l��Wн��剛��8�G�HIӕ�Ӟ�솲�CZ�~v�t�*^%҄��s�4���c3��l��K[�`����I�����afgLQ�ҍ����5l+p�����B%��V�4�V��F�4�q�6M�t�+��O�6Oy^Vu����H6Y�D��������9ˤt>�y���b�A�i����2��|ד��m�{��o��ȼ�F&-%�u�9���:y�����h�o�ø���G�$�[V�ҲR��!&�Sh�\P��Bֹ���pB��3m/?�b��j����v�T�t��E��Dt}��5�7��i��}'�y�J����G��p<�'�<����QL�i�cn#���������[��FF!L�	\�>snv"��=5J^�L���&-�.��d��	"BP\�J����X���={i�+�Gl���M��)x@��Fw\w�#��;�
�Ea��nޠ4�Mki[S;�����vGa��ۏ�.�N<W~��_��o�N��@
���,�Q�3أ[�{ȳ~�S/{m��K�b�A��r���N�)�-T���~��b���Ch^�;��;gyo\��祃�%�Q�#��'t����?�Ot���5��~�8b��,S>.���h�K���A�!�a�{��B�-����8�Q���-���K���u����a�vE*�9�8�69=T�YX�M��$���(�MT�K����⶚�/Q���k�ϒ3�Vmn�6L,����V ��G�}·|FtmZ��V�ڋ?����aS��l��3�ڟ���0����*_�_-�r������ae-{�@*�mj���َ;�6�`!�ޛ�w�9a�Z�
���5+��Kf����yh�~����x	�	�L�FI�l>tt�?u���#?�lv�>2@B5��X�d%������Ѕ/�4� ��ɺ�{��:�	dD�W����~�9l��Iz�\���RqS�݇%���Yc,?;<�G ~Ч�:7yU�?_: _b���cM�^���M�!}~�='4���9��o�U��3G�W�C��T$Da<G�˰�z�:E�<^䨬����K��'��#�.pE{$.%�m1	�6��K3x�i��{�$ܡ��)f�o����GzH0>���.��xm��p2f�"� %�ڑ��`�CI���w���˟�I{���1�J��aP�K��m�+LA���l�ڠ�:��}��Ԙ�����ɬ�V�7�r�d#_Q1�I��E���(~�91�AS�u���[����#L��A��-�%�f�������{�-,؜N+����[L�1v���O_���|/��W��.=�ڡ�#�m���@U���Fm�o�d�*��\�UV~�������،�j�n�?W�K����59E�/�6�tt�iQ�1���'��<��`-}���Kb#y&Y�k�b��oY|����#s�_�k�	iVI?u//�ne�4M�
h���SCp
�ĩ�Jl�0��j|'1� ��E��B����U��!��S�B$Z��&�v�w�a��i�.�Mpt�%M>�w��bW���Td �d#���Ϣ��mc�%�	$#G�go)��}��1hm����Ԟ������YvŽ�8M��6�RY�� ��9��&<WsK��d�Y8&|G��5脋���_�/���:Zr,�f�&���y|�$��1@�O��ɤ?	7�[v�i���]%��)�-=�})�U�_ޣ�on~�H%y�Q
��l���ʅ��&uM�����������wRq�bZM3�ts�����ł�[�(p�Kucec��O�+$fg,K.�)���,�b�7���Q��7��t*�ו�s.'��zj�9����s��|���_��r��h�G�E����=/���qN�P�*���!'��!KY=k.N�����>im�+������<q�̇��@7�O����b����@ ���-���FP��![Gk>2���G�+Qf���p;}����ڋ�z�_y\�37�e-��+/��A�)Ӣ�������~8��|�m�{@�츑���`��p��hEv����µ9�SP�6^ar��q�}t�C]^^�n���QLD��_W��^���:*ʬ��<'WO/.f�(�N���� ��ك˩�_��vFG?�2N���y~ �K��ؔV�7���x߶$W��b<W�����:Z�Z�ڔ�9����:�>���3- N�'�W�E�)@������*X -f,`*�����4I\1�%�F�*D�Z)޽+���/��7mJ�͙;��Ԯ����QߚHLk��2B�����jW-o���x���)ۆv|�9C�e"���D��[ 9��y�<r�>��y�FP���}~Ӛ�_���Y�M��/u�f"�ڮ��	�����"MR�����t�D�SS�! \���N���h<q���n8sd.��(��Q�M��g1)_���]��r��!�\�
�]h����h����+�usKK��!��������Q����v��ŭ�Y�b�L���@���%έ��v�X-_z	�ӥ����Zwnu3��+ �N_?*�2[��Bu\��Yo����(	;��B��q$@ hY���׻��(�5WY��`0ڱ�l���PD�x�v���N�{0�d,F����/����b5&���T�DFE�!a�)�"u�{��6�ux��!%2{vi�
i�����2E�t�Zo(w��j-����w��Ķ6�b�W��ԟ�60E64-�Tef��^���c-J'r�0�rz�� 슠 ����2�c��,�
ob��`����E�u��BXS�f(U⎏7��s�c�����Pfs`W�Oe��Z��	��FU؃��v˜*~bZ����'ح�j�f��&~�lP|�8��N��}:FϿ�ng4�I��#ڛ��b|��"������p�`Pl�̻��Am��H>En�����������+���4P�˻�TI�y����=����"���<���-����U�M�Jq�s���-΀��J!�(u��d��u65�;`�������b�
�j��Y�o+]ʮP���p!��R�ւ�_�E ��q��D�~��^�8I<`�{#5$7�LZ%�����Zڔ��/0s�OfUE�G]/H6B#�T�;��}��&�i��g�O#d����-�P��6����[��o@>�w����L�3����Z
�H�"UE3��yT1��q!;�����V�)�iKa� _�g[Bn�J*Ȳ�No�z�����i͇	N��uŌ�T0:��ίQ���}��e+��/ H_b00�y�µ᎖R!�����y�!i��ᜮ��]��&�f&��'|=�o;��[���v!Dd5 �ٖ̍����[�U���:6���"|�Y��W>�ׯ�9��u���---v��%`���|��6�y³:eXR��3���)����I�����z�R��'�	_ngy��S�"UȤ�<��1��g���R��Z�����l��Ͽ��I���^��C�Kbkn����\��1��G ��S�Vއ8�� �:��V�c�#H�F,��<�c�q;`+VY��_�ZĲ��n�SӏY��8����5%��9�E�Z|�͕�:\����/�׏G"
�`Bt�i�鍡o+�Ņ{�O��< �KC``����=�s�C�^��b�o��'��պU͉��?����lY��M�Wٝ��v7J7�"ϒ���y�q/4X���v�`�#Ho�Ǳ$���Q�D���4{r�Fʗ�S��%i�z(M���Nk����ё�����/FGA	%9H�� -��G J�+;='`�U�<�+���?Y��2`��x��}F��t��o�#�1�a��6X���2��}|�99�B���᪼�r�.�e�*7�ׂ,��n�՛�����Č���;Mz��Jk�h����_t"k�<�+�
�[�8��o�HWjƮ���֟�����_#��s��ksD� \SG�>��������e;��<��@�8��8�<#^�Q��M��G�V��I����ނ'��5������v�'{�����|�/�[Q�����������Yv�̞={@@�y�)HT�c�J�� )��L"��\���x�IM>��������6�o��o������L��:؎o�?�M�@�y�B�����d�cH��_Ǘq�����1_�pZ�
`���w�>���;J��7�Ҭ�2��������A�����S-|B�/yb[?�<m�U��Y��'�r��1��?{_���m��Ό�]��e�.��4�GSrx'���'�v�x%�mËN ���?~2�5�������X��y�!*�٣���b[M��ｿH$h�%�m~��?�J|���k��yNr	�Q�����>BS?�ÂǰG��T��g�~Z;(��A��:��B�c�V��uID��W��yp�yO���ڦ�4�1��W����խJ�抔?�	(E��L�g<sVP)�D��S�r;�ؾe�����g�5�Y�V�9�egGQ�>5z�Ay��HT�QW�j��<$�E���"5?=;p��ݔ�"��%���\J/�����_�h?Bs����
M�Xoſ4�ѝ�Ӝ��ڪ9J+����_�jg..砬�~gi����<O�����x�������X�\�
j6�V������,�K�9=�Y)ѽ���W .3���RV�s�41�w�1�0E�x�?������t�y`�h�t%{�������~��~P!o(������Y�ҜPR� ]������_I�X�q��Q@2'������?�2���R�P�}�c���NN�ْs8���ׯ.,������v�ќ7�N2��M?@�?���&H	�,��٠�*X.��U�	���		��\��&�����,��(�Z��m
��f��P�d��{avRC>}�劋��`�;�o��%@�@�=�v�=�_?��k����E31���%��/��J7Pm���5��2rY��|!H�����kU?=��u�gfLүa�\EC:́�d��*i7-�Q�_��=+j�Qj�*+�e�M����M��	�A��y�g�k��@�k��~ D�(K��KL'�EX�"�;#��QC+��q���c�J z��}���w|����. *��U�?�S+���m�� �a���� ��,��=�� i�έ75睮�C��[��/Q���LOO���h��:��b��	���c�� 5�g�5�5��g��]�淐G�)�gg>]f��e�)8��1�O��PnL��:�l���5<����]���l�G��=��pe�ha��~��<��`$
��F��c�6�?��@�#@��5�Qg^��B���7����9�Gp�q���߭#i*I��͜W��4K}�Ӭ�e�#jw�L�����s?
��$b�#bWڭ��l�l�����Ȣ��|$�r`�2ͿBЭʚ]J,�Y�zM3ѿ?ބ�D.�&��wi���h�.o�/v��+;ލ(�N���X��R�t՚�ݨS�Y紜�������E�[U]�>��(]zn������ Hy=����=�(��Km@�)~����B  ��M������hdd�TFz�� }o2
���w Nbn�T�2-���mC����;rHJ�����+%�	�2}��<i�`��C�t�7��\O������+���d;�?�N@��	%vӿ?�l A�i���^Te���wә}���^�{E��$q߳$<���A�'��n����� ����|kо�J>z�ݛ����V�$�A�҇�ӹ�:-k��<�� ����힍S�;o��7})M�J��5�v��'�k���4���' |Ŷ����wV���e����&J9�z:W���3|B!C��%W�����c~!��x����LD�8ڀ��H�B} y�Z�~S�L���T��� =-Aa{
|��M�ԕ���B���~�Y2�H��O�� ��4��a O��S�v+E�i!�����Oy�����{�����l��*%�K%�Hs2���;jÇ#z��3�5}9� =�S����Ԙq�wB��e6����b
�`�?�ޘO	m�3B�1�@�+��rr�W�;#1�8�:H	W%9V+֪]'�@�o�mЊ����e�� t�+���9�NɎt�ջ\29��v��#�r���3�vÚB�c�#(���>:����yU� �(�VVVY��(�S�D-�ۆ� ��G �e�;�(PQ�hS�f��K>P[ŕzaS���%]3�L�?�%�b3j`�X	G[���0�w #n{^�_B�s�� �x�aWJ��c6���.�C��v(�(+L�qx�h�đk%�v�|�
�A"�k8���ޱ�oV%ܔͳ�ې�Aw��(deg7B�\���ux
^����i&50-.@�쮌��JM�
'x�n�򾯡�|�v�,Y�6����3�Z2����:����FA��H@W�8i��a&u��^xjJ	4��ehV3R`��&�{V�فʞS�2�
e��E��%Y^̩�d[�-��%u�ē	�}}���&�t�y#p5������`=6E��$���x��	b�O���6�{�=��M<��ˏ�a���_���6��"��
�BB�'�j�*��i��cD��_T$��U��c&��`�*�Fo�7�Y��|3MN'Y��������P����prys�	�8��Խ�QP�ޯ�rs��yقz��oP����G�1��yݶ$����M�J��+~�������#1~�KS��/�98RC�6�;� �=w�TY|'���H8>-�]��v���RЈ��4�hQ�%���]�s7z�����cy�`b�i�p,]�pA����l�D�aVN2��`�M)�>n����;,ymF�\�,��10�@W1��zJ-q�)���ݙ�߬�h�Av4����Eԃ�o�!����SL�\��ls��UCο��l_^�~�l�8؆W�}���� T�y���u�)�`���6?<�)������ �ٻ=��3;�7@�����eu��Ln�'qOz�DC��+��+>w��E�,>���O�*L�{wz��P@�P<��"�&R[��q���uAB/�:!W���wc��6[�ڐ�XT���֌��$����/C�]�v���hhcA�G�)H)V)��kщ?$�"T�H�#�����3\>�+;�����^�-��7V{aTe*WL�n�ڃ^��_&ڲ���t�&� 9!�3W�zo
�����/��'yȘ�1�Ml_ll,?�����7�ӊ������i���f��~G�/���j��JC ��N�F���B7�c�E�E9^���O�JT*����n*��؜Au2���e֢aɏQ�^�jv�z.@��)@E���NUG�C�HgN��ʈ�3�3�}7�[����A�Y��{|��̍Y?~��W��	��}G �~�J֖���W�<U�4�8AR���� �/ ��Z��t�͈?֚c��K��2)��~N�r�pQQ��+�^^s��_�dK���6竏���iNֽP��ۆ!M�4�d�5�]t���B+b��������۫i/LHi��Q�{���ǡ$��U�Q�)��C��c��ߦ�b���G���9���㍔��-}2i���,��9�#�n�(cM�=�A�\bkq�	�[��)vu��b�=GB]�����>\3���'�Q�!��)k70'���(ȹtg��bpd�'�j���v�V�M��䅵;�rw7�g+"c}��N.�B^&�%L�\]IFKE��OL�um�Յ��4�H��?G�Z�c+�ut���[�*�u{�~sۚ����_���t&>���kj�#yS��>}.V�}�
��V�Ì�u�eA��V��e��'��|�/68$�^�R��d�oꯉ�}�iW�C�-w=�ܪd_c��kf	n��3w���VM�sz:�����-�X�W�Љ|_qMs��_?pU���	O�_����rGv�jQ��z�� Q��xu�k��5����W+��W��y��/ζ�Sgeee��*���|�J	���6]:����5ve���E���p/~����KGKK�]���@��3U�/_��
��|��Y��o=�ٝx�|n�p�R�ѧD��݃¶���	4�MW;l�col�!{@qqq�����JT�Z<]�ݟlv�J�4��0�ӊ&)%E�ű�h���x�X����S��x�l�/О�6�C�X;x\Kp��<�zE>���Cb!�m������ !��o	�M�:�'�~�����������M�>}
B�;B���OG��o�{��ӵ��d�˰}�O�z aF�豮��%I�k|���^H�����!d�!T�ԮE�g���z�����Ż$t��h��њ(!14<��s��"��R�Q%�ߝm2_��p��w�ށ���<�`No&w�����)|�wX�q����$b��߭�1k}i@���hvj�kË����X��yLVS�#��$��W��Т{jġ=��׏��K���@��,v�UC�jj"�/�H!G��!i)7g[���&�HK�Ĵ=<<���]�`	��Xt��G�T6����m1�;�z,���v!��%_���k�Y�Nݥ�T�����3-)l�d��B�VW�kdi�;99A����V�W= "i]t�|��g��
%⪼�� 'C�j����/�f��o�10��w��h
���J���3p+�����+�K�#"�R卺�Ɂ)O�[V��O
���TS�ᆃ���L|3�����2������Z`1#�(@�Qv�+�sg�N�u��ٺ�����UA$#��RU�ɾU��Ew�>��&��C�h&�
Ʒs�����Yd;]��˃�h#BJQQq�Mן��ُgyF�������n@=��w�\��ǩ����O7$�;/@�*R��9���c�M{�$� �&�vp@^�d��ONNf���ԟ����0=@�m/��$BSиM�딦*����n�@ۣ�k�r�t9�%95�ֿ�2�#�����x�~东�l�7iI~�ؑ����s��I�����ј�X���Q����f����˧�_D\l� ���?�'��RXTE4��R˕����Ȳ_FMM�=Z��?�gj4|�o`����$tKIl���H�م?qT SH�<W�	 ��URd@��e�Q80�]�{�R��Z�.��b��S���C��] 5e��������w�r*e988������*��E1�e@2
��
*�s�DE@� A�E$I�X�JQ� X( YA$�R	*I$IF����t�s��9��ޟs�{�j��&3�����1�Z�/�h�S����;ݥ�%iHt�����Ne��G W�!WD71[C�iU55 ���R�֦^��Y�{͌���{BL�;�|���x�n��76�
�u�x�]^r����M�m�/�'���]�-8h��|��(�7�	Pd��5��O��qAB}�O�C2J:�"5x��A��`pS���ն�����
p�}d��hN�l���ȕ�u�_���Uf���v�up��ŎBo��))���C���"P��G���a��P����N�ԕ�����]�/ $���Pf�~�Ǉ�jj�?vm�����{9)�������p�R��/���6
�±�h���|��p l[:�����(Yߨĳ�7��g�����ff�,��i�	�o�wE{M7�J1�����Vq��Jiizn���{_^\z��h���,�0��5�*�NF�����n*q�`�Y!�+����'J·<��yݽ{�|�5�gֹ@�� �h��.Nj��-:�iu	�4��ÇU*�K=P��7�XI�'J"��7:��7��q��@I@�b�#Q��b̞����,���o\ؘnF���a����; yV��ǡ��	�g^\%����?��m�����F�ۛ[���w�!��D�%���O4��C)+((׻��i@� NMj]�K[y�N0{X��Ā��l���6L����l$�h���!�jOq�B���_���a��ڐz����=�	�k	
�Apz<r)�Z�vOy{��������P\T!�̶�����}���7�RJ9tu.���Dy�6A���t�p�N���ӟ��:z����������uTJ�4��2Z�/�N��%]Ȉ�X/yɩ��?F�q�raP,� ��(����]^�}�nb�7k��i>?~�Bsf�ʡ�rʻ
�֬.��͓࡝��,vd���0(���֬a>�t�<	rQ}����b-Nr�Z��9u�9����6�B�t/�!���<��� `�{�#]����]D�L���Ij*�Tu��/��t�y�g�B%����M6�^���* �;��L�����]���ڔb� gjC����u�&�nnn+�K�ښ먯�펽�utt��g��d��6�z�< 8��}	�hW+�2_��Ն��������v��}K��|��`��"��u�LϷd�����S��8
�B�;_U+����P8oC��p�?MKK�g�tV��<���ƫȗ��s�:�Jr<a*����{l�եw��D{�in3_;F��%��mv��j+:-t藽��Oq�o�P���u�ߠT\IP�ם{Iq���~­�3�z��nQ.jβ1h�uR>��{�~���	h����?���x�p	ڬ��mg֧��(�(������4�Tܞp��՗�{��:�{LX�Lo��������EU�><�s|ݷ����/G;I�ػv2�y��U�꺪��0�X7��ʚ��� �~��.��z���
��S
"���N����/*���V��ԟ#�|}g =�v��[h��l�N��3_{����(�TVr�0J��%��� ���|7�>͑�m �bߟ=f	�-:bj�k&�	

B��:٥gN�����������ݭm����`�_܂P7\��AGL���]]t�z�g�9��	,��(��<v�~,��jӗ�"}[[�� 9��赆���~�a�K6C���kٚ�H���A��4Y)�I��j�N��N�B4!ޝ2LIL�<�bl�\�R�P�N�������l��.hWp����Y�Ke�.�ԉg'��W�Q�, G]]B�y %o���Q� 1�.�\�+S�v���P*�C,��1�� Ud��)�n��9�L�L�2�?!.�Ƨ����;k]��O��$m�&3
v�T�i� c�[|}pN�%�����ggg��:Z�[��<�n�"z�H$�^X��er`�K�=�+�9�S�X�����%)�	ӋS{�������zܑ��<�2�� ���#�op�411A�+�G�窕Q�L�ϡA��M���90oA�������؉��X�QgRUJ�[t��܏FQd�.&&��5�;@F�?����������~�3���!UO�J�Em���$�䬔�^�a��;���٢��0�$��yg���~TYϏ����wBѮ9ˇF�o߾y0
�G�����	��p	 K4������߫>����(�/vbA�5]m��p~MCd�ʕ�[v�n���ă�`9�;>A)I��^,p�������9)%�(��o\�ˆ��7(��-\|(6�ڡ���Hɗ��15i��@�b_�/�]�L��1ӓ�0��~~����T��h��"�P�������*�ċ��VS��N>�S�c��w�b�QJ�ph��@ݾ�0p[��&����̇�F����/�όw�?��#C@u�[��{'�e�bR�)�-a�"�O��?��z�}k�CCf�~<��,��FH4�Ywȝ�؁36 ��}ū����]��n�?݉���(q�/���N�}��sx�]�9�������KÝ�.�~��k� �]s� �Q�0��E"����)1qq��欗-ٙ�n}���<���~|��>=�rs~��Q�f��^m�366��ڢ�:Z4=h���ޟJ����ڲ-��	`,亮��h���;MaKs]��mTV�(�]UQ�:/�ܦZz�u�H��8 ������W�v�(!p�ݻw��س���nq�V���@E�{J���4��	7�^>�%(%F����-���o�������xqq1�f⿽����|Z"]���'R<v#$ ���a@��a�@��H�)���'�ԙ�~��;��Hî�~.��FI�
=eA��g���F{�I���������2I�\��⑰�nY�0��S����=K��!����;���_N�8���+f�]�ho�vA /?8]Hq��y�Y�'��6g�@�'�/t�)J��l�~S%�tDT$�l��$����˖��b;F \�[^�07�2����u��s��},&xk�N�?;?E��Ժp�iz� ė�ci���$�<��Z[�iU��]�v��O�갧��C~��"��b�ڊHii�֎��ٳ^��[Z�RAA�oOn�|��N)ccc� ��a���}_��,����֦����k�P���l}r	�D�_�h���S"���fH{*� +*)�(++���馶�:���S!��pG�J42�����ɨ�>����#��"'	@lA07�4z>�B���0���ͮ]?jʋ���?�M����S����h'��+>�_M5Y	O�sjjt��U��.dX��
EO���v*I�&�H-.{���n�0A�Pq�������ʵO6�d�n���.�X�Ag��r�4�N���|�ɴ6x�{�c��f#�Y����I�ZI����ж:��|�;���^D�oș���u��6&��7��GBhE��a��ND����Fl��c��X.��?��:��_x}��0��_vTJ/�B���?
�Wd��ty4'!9yH,/�Q__�;������1��8q��?	�E�rt۠��+�.���Ru!`�Ƒ��ne=�=۶m�\Z��k��]7��8K1Kq]�b�/�E�C?&��#)��)��W��	)��`�����{�4��0Q��![dِz��U��R�����A�)�.F�qU��܉f���6�Ag+DZ�h,:����VԺ8L6�����_�n
	-�G�쵒cx����\gz��/�b�dz�p���0�oW�&���!,�<�I�12�O�B=���I9�/���SYC��m����&`X��J�>ϥ�9��ո,�ڨ�Ol�(�Ӄ���{R��7����8��kmà��68r,���Q���i��\��{0�:��䯓�N�:��䯓�N�:����ѓ�{��6��ݺ4��5��ţ�����t��c���������U�?w����͜�k�^��
����y�ê���_��o�o�p��N�[��V�~�����Ͻ����E���_	�%�����KJJJ�Vɭ�����X����(����N����&��������c�S�Ɩ�TTjW��ڸ�������I�N��&�n11�S>�md�uq���V�'M�V�'"���4uf �֟�YU3�u��~�����=�𵙡y?��>Ӯ���8��a��$մ��.�W�B��<�]\0�7��QO5j��knnn�.��Mz�`�}���ƟW�)k�H���&¼:�/T�:�pqq�V�2��l��ѝQ�UkP\�~]����8��:���TƂet�X�O���ǻV'X��c�=���b�����Ɣ����ʿ��K�/����8b1Iq�2�i!����Aܽ����$''����E�s����p�]eSS�e�����):F������!y�W3��{z�'���Pp�E3�;Mn�֞�MV���jZ�FT��@�0��������K E˭�w�ۅ��K��E�+[w�ۺ��e�F��[�:�L���ެ���?J�_	�%��_	�%��_	�?!�q,��zX�veeҽ���xh�'Iifվ�ȴ�cV:�?��N��8>�ƭ����O���s�*��_l#�o~A�?����K�/����K��;�$�<�R���9B��<?��˺���{�2>*h�c�;q�С#��B�_����]�_'��u���_'����I��vJ��#�9}P�l��s�N�|�^���������C�ˊ:��;���x�./|Q�n���N�U+��>��5M�z��bk|q���d�5�|�r�!�耧�����3��e(<e����Q�M�چ�s�Tda����!�%�{�8�K�֜yk��a!KA6����y���{��pݓ�X�G��T�y�g��"��):���z�z,~�GXNz�^=>n��vk<~	�+������b�y�ؙ8�Pۜ�3d-?}�:\�c�J�=p_��$���&""�L�JL^8����JZ�����ԑT�_3��Sxn���n+��D�����%8��R�ނ���r�@�
8�"��󔽐�n�\B���k��QG�c��_-����t�*"2R>_8��y�8����l�D��3��r����)��Z@!��U�i����ИCX/��`]�\XT� �=nx�U�9�#Ұ���a�Ǯ�Os?Wk�2Mk����7�S�����Ĥ��`��8f���s5
�)������8�,��o�n�#�ʡ��)��A{��o��֒7����Hx�3 E��k�j�CDr���ԏx<]�����H:E���oOi|�P����j�t47:���* ZD�\��QL��'�s�G����}_0*T?��H�El�!�`���[G�絉��tqr:��Ĉ��rK7e١���Oc-X��߮��!;E�l� \�_@�*�~&��ؼ������y����������J1

W�j�&���1qV�&�Fq9s��YZ����! ���U���-�3����_NV��l� .��dl�	��C�����tOn��A�B�Cb���2����#�����(����1��j�����+zm�4�&��ﭳ����!�]+B�"��_JRO �+�ayO(x�I�qe�9��a� sH:8�ow���h�y���j���\Ľ����1q����p	8ڢtA�9�$g���Q��v����D��L	��$A�h9/b�Qe<R�_k��	���v��}mNN+�H>��#I�f�I��b�wY�an���'w�"]�����r����?���sZ��:ϓ#�c�CV`ĜP�EƲ�^sZ�c?��i/l1g@�2�@8�g�	1���r2�b�!/u�r���p�u;���l%XQG��V�`�O���
�Ӓp�_���H����(�M���<�7Hr!���T����ɍw��z�p�_�v��,��>���p�����]��Z��_�E��q�UQ���Q�d.�G.�R06[�& +ޮw���,h ļ�)f�M\�u�q�Ć7� 5����2�"�쟝���7������!��f���,���S|x18C.���^TP%�S��8���,�F���w�<r�>��n9��J�Һ�bǑ��U|�!RL/ɉ����?Kv�(��9gD�j#.����,��i69-������X:�����x�w�������3��d���Zةù��,��(�K�vb�
ƅ��Ew�B�w:)ƪ�S!��,�q~z/���[[li�
6��0�zF�e|�Yh��B�6X��	j_8�L/WUp��v��е
ӂ���R�/�a�C�� <����gh�'.Ml�_����cd�m׸�J���l.��Nx��{6��. !�q�0|^�7Y����_'�\����Ts N|j�;�g�*%b�F�r�Z�KG�
���:�����.�
fB�����뢀�O:)��B?��bH�:�zV�̂�ܿ�q2{aԃ�U����+t�[���L�UV۟���8ƿ�J�i(F������ �%��WYp��m����a\sz�Z���^h&_\0�OF�t�@{
��	V�lbG��N��r����&����>�[�8Ym����b�?�ܽ4^�oGvy� �P��, �w�A��B^~���귰������Vy��<[��A�8J�*QӜȃ�������&g�"Ռɇ�OY៑���wf��'��ħ��$��〒����C쾝�r��j�������	�V~Аm
뺩������L�h�`c~t��t�w�3�M��>��V��8��cϥ�J�&���"������s �L7`��r���9��BAz�����~���y_`�>���M�`�1�ǉ��=�g%ͼ�P/�%(y����6��6ui�+K? 8O��7.�h���D�ry�Q�M-�zvo�M�L�y?� �cIc�b7��Ә��;@o/,X��y���Xd�qb���6ֶÔ�O �<��<}��%�7�fi�-��`��ͅ)O7XؽUؠ��\A������`�����a���s�R=�%>⛯�'���|g��H�ЫM/4�K\���\��W�}�I��>9���֦�ʣ���6���w� ��љ����k,����*��p�aFP�M�g�x��6�]DPO|=� 4f�:ݦA��u3����#,8���&��Rk�!R�V����=b���rWS�sL���J����A$X��y)&��~��������O��`K��j&&�����;�S���F`����DԼ�6�q���r}p��+�{dd rY�0�j�J���αm�c���Im��l
���!�:�g��%�7N�����L|f�1��N��z�+`;���������TCқ�0�Zd跡z�k�q
y`���i�X}>I7䔥�o�'�kz�Đ;�pݥ��(h�5=,������G7��Ɔ�c��Y�ۗ|]Km�7�k임�@��#�+�u������áa�K����@�G���H��Øh�=M�!���U�]�e�O|m�N��#��q���:���]a�5�Bhk@�e��@T+{�eh@�)��;�h{��'HM�ml���h9*6�z����S&����!�#1	�v���
��	�ȸ@��a+	�w����i�҈�ݗ�m��'fx��>�A�YY������v⵨�*�w��0�D+�Zr	���6٢Q�C��M6!R6��d~d.N;Z���e��\�s�YμfW�qW
�\>�����.���� �?�u����,�CO�+��ǧ�!4nm��pn�5��n&��/�;P�΁l��p��d�h�6�"�J���W@�R}*oB�,ݔK(3�}`���{�bsV��c���(�}��'�[�Ÿ�}��OQόb��Ȳ�b��e���a�Ox����C�hހ=�	�&��.F�@C �a�=��xp����'ۇ�������δ�|��7�6���0Қ��d�>����)��Oq!��D��,��k�B���rH�z�6��F7QE���d�À�BP����o��.��pֱN/�G��<�H� sK,��F7C^P�	���A!-'�;�Z"��� ��l��Bl��]��˴R������e���K#r�5�̸�������3����i�Z%�.�ݼ�߄���(z�ly�~֟}OT9��.�ԯ��G�f�r�&�hhvS5q~��s��n�X����(��K;��B3"��VD-2���"6݊ޮ���Sn���� 0,a!���������\�M@��+]_>����0�?��u(I� '�%�e�6w6�;V&4�	��";�__��u�)���_i��P�j���|nf����n�g���^�h��.���t$`���7���A-XmgIo��|�`�Nm���Ǟ':j��]���_s���*+��Jn�Q_�t�K}V�{���<�)�+8<��f��@^��@�|6�ЬCF�r�]�
��j>��р��֢艭!1Ff]���Z�0�z�?�tJ.��;@.짉����O�]{kA��J:�g=�u�\���k@G6⊯_/i%%�+<���b�#�Sh�	��ݏ�����lA�3D����~�j���RP�VH�d�<�����I�%
L����w��}�n_n?ǂ�z���+��ep����Y�S��R-j�_ތ�� ����3g��W���SX�˚�C�B�*�4D�pV�8C��{�޽{�/M(r��Al�G�[�\��.>#]+$:u3�'.5h_�"5���Ėk��vC%:>�r��v�f���'�>C�B�nW1ҙ��E<�����mL��pt����%0��)Ȯ��_M�q,Ԕ�a߲/�{i`�V]~�~����ǘR�A�p�3eB�8hܤ V��1�
C�1��ZI��WZX�>�'!i�*�<�C$����cx��#�YO _�;Ԫ/��� �Mk��{���@�n9r�0	�?��Ğ:��n�S�2�5���KƅqN���N��f#r�gwȸ��l6������!.�g��2������ܰb�*8����E���2{˛mV����{��Q��6���O�f�;�3̗��D�|�l�������N�ޕс"�	մ��$��Su�������(�W�7�o|�}(�3X��Dmt�Nb�q'-J�+΋�͞�U�����2*?�9�,q!�"�i��J)=y�-�Wi�?�ITWX�6r/a��.:���k��
Gq��k�r�uM��?�B������y0�����@�-IP��W*�}*�ȹ��!o�/��{�¯�X�����M� �S��
u����"���R,�R��0�]��;6���2���5Z��jy�g��e�ol���n��ij�� 1\�N��CF�o��>#�֣���,d<Q��	�IN�Ѷ ��~[x�6��yiݯ���rd��ŵ`x�]����*�����؆&�"��:����,��9� ~�G��������S�T�D_R"��k�$�両�Q\~��e<�Ϥ@|�A>�	)�,��5��g2�~*�I���D�瞫���j�V���������>9ՍR��߰��%��ʎ���02�C�����Mُ��ߡ��ˢ��΁��wq��I-�n�d�Wa�69��	D����-K�����E��q��Ap�<����f�S��W?C��~���~*�< ��	�6����� r���*8#����=N�t�*g��a�N���A���e=l�}�y��CW �m��yn�]���UM�OQ*&9�ǿ�q��Cv7�}W��,c�I"
����X�h��e��ot�ّ=�u[_5�`�B�����V:T��!��D��"w
��� �tr?����--�B�����1��{����d*�=�dԸ���HZrG�:�m�BJTI�nҾe��KȺ/:W���'�;Lv� L:��_�����n�����l�^&xe&=g�&-N� ���G	Lx6���T������ƵB}��-[���"�����+��\J��"�l jd�uS�_�X�cu��d���A��d�c����fA�Da2���'�r�5���8�\f��{yXY���= Z�~Xy[�5Se�Ĥ��o�P�.7���~�lHe�b�i���c|�ktg�>zzŸ����V҆k�O�'���^-s�ƽX9�#�l�*�[����Υ��

fl��
�Ė�?�/�����=�#6�wkY5'4�Ҷ��%��5���:�鞁r�& �q499?�:M:�q��"jJb"��1��EF�J�r���|��ŀ��'1�<-�w��؜2q�iO�4K������c���w[�ǘ�C�V@:���9_"��Ecc״����bK��������[���z_]�͗�l7���<�{�� �w�ǌ't`�i�r1�ѳa�l'׊qI�s�MI-d��12�,�u�=Ed��ђi�͸pq��b�����<F�����g%ŵ��O��?�A�u���~2I���V�h���G�c�k����N&��:�X6���s��@��A�bF�����cn����!�H���'�D�g��`}ExF�����nKI�"�FFݴ�3D���3�:}0�b�z�)Q�j�֍���ñkC���^i�
�ǰ�A��2Ϝ-��]�Q{�r�Sd��iG���n��OC��^7D6�Z��5ӄ�}͊w����ry�K�T������;�xVJ}�ll��8�O\�L�w���A{�+�H{fjP�;�+�$?w���>j%&%�*Ӓ���%�u������f�5a�շm��@�H�xll̻`9I�t����U����k��M�'�u�o��!�do��[)�W̽ON�\�15=��B�U�f�3�#u�L�
�z>nQO�B�=�>��M`h�-�5����ѿ\R�}1*����W��~zE��ӥ����E��-��y��m�v���:������;Z3���?>nD��]#��
ȩ���&����,xz$q�K�gO�E�h/��>R��l��:9��4u�191���{��������i|�9;����M�p�Zq��n`�J��+�q���*�e�l�ciJKKc���,#X=�Ӳ�!p�����'��Ƚ[�S�J���-�M�/�#X0�z��3M���L�5���$�Ϛ=ֆ�|z<o4��D��F>�LIV}�NTd��ǉ�B��L��6�H���]��M���㉿r0�;�]�"77��="��T:76�FyMLL����z���=���0n�B,EKG�O1֦cx�삠�����qvn.��2�%������g5�J�E�ʑ��i?&�=�o�6p�
�J`�������B6�.���c�����BB�Y�sXM��w�Qr�&���	��/M|C��MУJ�UeG��MN��]~'<���b���."0y��z���\�i_ff>BF_d��켶��fnn�>Q?�s�p{>���� G4��+Z�CR`L�v�4(���.�c��kkk��O�'����!M��kzu�91���bbb�q�#��*������ V䬦����N�!.��7D\@���2��I�N.�8�9U�	q�����t��e��\� �llƗ!���[���ϟUUDFՒ����7�r�1���{�����?T8�l�ZPw����Y8/:��n����ߡ�����&FF�ꞕ������ �= ,�&���%�A�˱�x㨘�8�|�E�$S�P�M}c��=����\�!��v&ϊ�����+'�^�\�¥�O��и1�+d�Ut�<���׸�Є�_м�2�^�(ڟ���-@�K~�5 �FH<����3����-��0���CLE��9}�\T��S�h�B����|BBB�bbD*&��(7��f������]7޴���Lk ��w���@���Ї�� K%��,����I4���Fsv�
;���N{ǯoo�u寨IܐX�~�}[fN�6WAP[s�D��Pi8z#�9'n_�o�~{��s���N��!�����RKG���@כ��e����>��K#6�4�ie�$����`_�'2y��/���^�y;{���͛7�a�;W�|�G���P��>/*n[��
��m/ �s�a+j�.�"�N��ǡ���Ӫ�[3S��cj�B����1F\�tsEVrH�]���1>ԍ�^Ou]]@�����[��åpOP4))�o����pT��i���~����`SSӨ6+��y���ݵ��|{s�r��( k'"	<�Dm�O@��БU�Mΐ���u} �ein~�'�T¦�J]�4��t�~��h�� �V��3�ǻx0X,�G����"��H�.�q�CF�y,��Àx[�?�c��>r233��Y������J$��0�X�]�(�Y�S2�0 t#0���V�%���E�4n�E�2����T���G�#5�Ͼ��?��'��TdT]���`���1�QD������
�Z�X��]M�2H���J�T�킮z~LD
��M����5��-e���^;d�mr�ɿ�.��JzU�B���ԼCJ���˿��p���]-P%�@+��]�9G���-C��%?)�(�"�nH�LY�g/~��wO��Y0�Ov{��{�/Ϲp��WC�ys:���:�mU��`���#G����7:PW�����?r����Ȋ�Ө��M�Ccݥ�[�5��| ��))(��u�Ƙ����-�eX��f�{��$ҩ'�2��1��J�srj�����zj�%�U��r��=��޺���YM��D_!�K��;�N�<<��Zn]}}��50���HaRS[Pԩ�q_��h�egow�ؒe�ae5"I��I������)��f�Aitv2L)g��ډ����}�o��"��u��1���$!�y�$�G��H���b�5S�]Y�M�íM�۷Gx{�nB[
�n�C�j���P�-��~�Cļ� 	���Mh#���[������ܹ��z	��Һ��M>��eVf2	[<@�Wij<522��5��R�y��{�@�цJ����z�F�E�8��@���?�,=�0��7�d�/MmN��cjA/;����2�hqG��S���J��>z��/����[ ze�� y(6�5��C8ڇ|0��s+T���S�k��������"c��ivP�@�g�.���N�s�n��;Mr+n�w���Nv`��z�'�٭w�r|�?����E�1_���Obr�7[1����#�۷o���& B�!
bu'�Y�<�DCMm�]� �6�st,��4��7���Ä�L�V��x\hZ@���˗S[�=.Wmpշ7N�tS���8����ٝT����6m�PV�M����ַ>�t�hɞ��j@�P�U?z��ᄀ���pj 4lq�{i$��CN8#d��X���Kʴ����Y;bKS���Cj�m��)����H�K&��>��[@+P�KO���H>Kk�@�s����!���o]��X����i�jԱZ�xxأ�.�B�CNK���DM���}�o��N�&�����13^��P4���d��}呚k��Aew�2���T�]�X���Dj	��+s�i�Fv�ͷ0�(����ଔz���������(�7+U=wK��(��?["��J��W�/Í��:B����w")�AF;�5�����J�,^��>�Vݠ�&��:��&'�ڮ��ȓh�T�K7e��k����Ԇ�<�ڣb]Yg����e��n#Mŗ��ًuwN>����^5�#+��.�8�x/GK5�uڢ�iӜ8'�v���m��2��ʴ�Mk)H�4���S9�&����w0 V@��,o�T������,|����$���:6��P3557����K=���yAs�[��qԽ(����kji�����zpȱ���J��.��~1h'��E���`wW&鸰z�ƓVVFb2ci����"����������kz&��s�[ȵ7�~��e�w����^ʳ�>/��� �� �B���&�TTa1N2�	���
66�������ή*i��Lbaaq���N�mjBX��~����Qp�YJ�}G��~�������xR����k���ׯ�y���"�yY�H';�L���2��L[988��z���/t�r�L#_�~���޲A���7�)�, �(�a��H��Xse췽�x �W�`�+��)�{{E���e�F}ikiYhyj�vȲ���7�t���j�&IpΔ]N �w�b�b\FZ�2)�_H�A��L��&�Z1��W	�-7>^P6x�FIz�G۫�/��VK|ЬGq$C��ec�z��v���
ɍ��Z rm�rRh�v�nm�M�h�˯�P�.�}(� PX���aڳNz����t�ŕ��2�
���?��2�Ҙ��^��2����j�;_t]c�Vbr�"�s��{��8:N�*��]E�[r�n!�9����"55n��ń��Yy�@陛��̚��g���,�����9�O�Bu.�C�Ά��I�$�I���z��6������n��D`HKD�.�� ����.�֩
���Ns�� ��V)�}{d
����tK�'[�k�x�+�4S[������*PN��w"�p�s�K1o�ۿ@����=�����Z�m6�����Y֝�7���E��L��ױuD���*h��>��અE� ��
4
����$�������h�g��Z�d$��u�'T���
l�Ҧ �ՑWs^n��cU�67��Ng�d!�L�5Ԑ(����<{="T̀D	wv�Ia�z�h⣃�1�p�*z��1G)�?al���8�F%�Ѵ��8���f�00�=�}�-""K=��+���k�xE>�G|���6�~��N�lh3�X�G�=mL�+B�l~��}��evv(�n�j�t����T,,,,���%�n���t�	1���7��X3g,�x94�Li�L� ہ���p��`6��L\F^�n�r�(	$�,p�jkh@M��ǘV6 ��\.L+;����4>��&�)�&�+Z���UUc�JO����6���l�� ��Dv�j�~��a`J׹�����?����~/�2��'j�M����Z��$5s��O��lc�4�!P�t�J���S���L@���h��a.�lZ��&��L�Z�88iXT�ӷ�E�S�p3��27�]����H�i(Jh���tV֝'����bL��:\:�L���w,�S���TTTȬ�"X)Q,{��0�
+�E�Z<���I��2�`J���o�t-�����P2?��i�U���"�0n�-)�![����� \��Ą]���M�6b�I�)4�n!U"��143;����XB��J�ejj��]`WK6�k_sች��WR��na2��#�#���0�5S��\�)��.S���a@ R9c��a�Q��`vww7L���\V��\���Yꠦ6���p�i?�ǎ7ͯ.���l�fں���J	�9�)|[Hi�����,�"��p ���e�(��?}���������2�00��I^��ؔ�W����WU��9!~օ�%Ւ���X"b �sT�����n�qw� �C
�k�ܜ�Dg�q0�d
���fT�Օi��u��)�*4���*p����� 3P\U��S$���6�J��a����S.�U���f��R� �.�����<g���^0��i���]��S�Z"��`)�B��d۠���D�*wF�#k����	� ih�2�7��MP�(=��F�a9�����TkI�7a^����f�Q��T �$��=��ʿ���m�����D���o ��q̏IèP��a�PM������=>�R��x���E���J�ؒX��\�2�M@�]pWq��2����Lʋ�O � HQ,��`i&=7�y˖-��f)�5.]r�K#�J�0v��r������W�hn�LII�#���55b&���->�����U#�0k~��+�Q$�uV���ٚX�+:��N��>gep#@y%$k�ǏgT�f�/@���9�@{́p�A�r��#j��j������x%%b[22������� ��%uu�Z�<�/d��c��DfZ�պ��-˿I/�j_:���JE��l���f*��t�����V��CϹ���=I�� �9ҌT���
h%���q�Tzf����3��5�o��7>��K�1�)82%(yN|���̀�ի��4J��]rJ�VCY�ꔔ�Ҭ�Ps���V�� �0zw>��=7�"��<e5�3u<Gr�a,������^~bDtG ;�?�829��R"�:��8fP�=Sc5������v@�]���K7��;����6�r��t����-\��0V�3@q�Z8<B��hqhhh��wS��m�N6<�[��Yz_�梁�_í�rҳU���%��ˬq�0�M~���Ĥ�S�=i��T0�N�ѻ�;������<�he� �����>1왮�eٜ��}�%*��o��%�aEg���x��T�P1��K����.dg��ڑ����.'��k�v�bM�o�Om1|�1��s���������R�3<����c�n�6d��I����Fl��JQPT,���|�3��s>���0�g�&o�4�h��秙p����d���X�����V0_Z�*����،��H�hA�D���΂���w��۾Yv9�˷�)2�8|�M8���.$�`g��Y�Lby����Υ&�����f�Xd��͎��ߟ���hLlF{�%T��a��1�_j��1u�c�ToqL���m�K��K6GY%Y?/��B�:-�;�y�^W��x��WeZeڢ�vxG�9�"�e0",��nT��5y��(��2LEؗ���QC��w%����1��O[,���Fs�M�S��j	���������F��[�����a��|����͛2-ڊ����؃^�$�.V��j��c��`A^̲C�㽕����������#��)������"@p���p�g��C{�2\O;}$�sN��d�d)#0���Z�?���RX��O'k=�ˇ�@RL���UKK�o]*�*�&��֥\*g�b��\�G؜����CK�T�C��:BRR,�}�'��u�j��'6��a��r�z��q�>ʂ����z��m���>���R�܋�|?�%QM�j�g�Z^�(+��㐿De�dZӗ/�����򳨑c2<����G#=.-�,��.�����@�e���VҲ43�?Y	C��"����mN��ab`�	��]��L���|I����Pؒ�����5]i&�Iꁵ9~��k���{|��^]C�Ǝ��J���>+�������)zyI�� -S�tN��L%n�����֝G�J��_љ�"��-����M�J�V�]֞��@�3�
f��I=9�?;��T��]d�1��(x�ºާ����U�N����R	Koa��3�L���Ց�����h�\����[i��ӳ��N���[̓���h�oh>���իW����M)��3���.d����R�"
�J��VV�ᄱ���|�������S��O>�:U�P�ѡ������#T_�����(��$��ob�� �Oc������p0(v�*�C>z ��S�-߄t-6�i�`f"Mp��&�,LU{E0B�#"��L���i�Z\S�g�3tr^QQ��"�!z]}pP����H��{��>�)0=kK씗�?�onn��͉�>�R߯�"��$,rW��)�.��R12�Yx[��o�fW�,�3�\R;L���4~�qgtt�ѣG��-�'|�2�������~___^A���ü��dӵА���E
���%��eZ��ӂ�ެ{������u���Ij;�C��s$F���5�7�,��$
n*bA�8W5��&'���rr�O�k�	j�DD�UOx��
&�UR@~Dx�T��JOW�����L�LYy�,���.��oE�����B�y����1	�a�J��/"�W�� c�{=���렄t�"ڎ�oǤ�i)~���0&�@�}������Rd�g3�Hi�Y����%��=?;{W��� UU����H����4������O�Y��e��{���U
�����VT"�&���&��h�����ՃW�ĸ�,�8���i@b+hWVY�?���:��Cg���������߿�cgy������5̣;gB�͹}�O�-4�i��7545�ה �ÏS5?;�Q����^7�5,���SO(*.>	Ѽm�L
�~c���f��B����k����>�lM'^P "ǥ�ӥk����D�s�	������8B@awτT�$;O"j�!nU�����*~E�4N�9� #6IUZY�j*jXu���Q4�f�b�ڈ�6�����Ϟ M#!!�Mz�4n�)b.#��LP2-�*�����5NI���rH8�2�wg��{ݐ���O�k"��s��J�N$�Tu��O���,p�9��GO�\�ؘ�职o�����s�;�kk^�sDn�dg7�v�O3O+�^\\��4rS+~�X��*.6���R.OWI��)�I���悮�/?ջU�?�,���֦TS�=C<o��뙹��W�?~�8U�*�N~#'�̮�IC]]�ʕ����g��]��J��5����Kt�F4O��@<�r����3�����1fM���>ȧV�,��SV;�ip;3�rB�>��%������Ԧ =(8X{�f��'��p�L�}��u���P:�f�QU���i3��S�)S	�7b�^F$���9iA�b�y�0�(����-�v��������m�?��������0�H���
��lS�MO7�ѣ4S�]� ��r��K��&A�x�t�޿iӦ #M`ZI�b�}����8<]��C��룁*�?-�!�Ѵ;��Ғ���/�¯߰ӥT��
�$ǝH��6f|R�}��eF��x@9$����L��c�v~�0 	�kKS9'���ܓ����{�!�8��һVݡPVQqP�6��! �U� ү����=�x�J���:6�8���
ŷw���aR�����ԚA���Ƕ$Eq��]��yKK���EEE�������������xq��	����MԲBBNk��v��D*R̈��W��ޙ����<�P^9�>���uu�ж�VR��+��	Dp�l r�[��)㌐h�_{�����\=�C���_����d%�C��!�:+G<��>�ߞj%�}{�s(;;;���ӓ����z�����ԡ&io+�'Y�������H������玄�C1#�� ��sr�ʍ�Q�#EћY8��ޗ��9T�ځk)�s�&D����8RU���U^VVXX(�9NP�O�1�755A�t��^���gv��wK�LrQ�Ӳ�����Х�6!{&�znn!l�����~H-?&��N�<����1I<�V~Ю=~��5J��s^k��F����j��vNR�����{�,'��e�ڇ���m_ߕ��@ٔ��ą_[%��|�u���ʍ ?���e��)�k��`e͕t��>] 1)��e``XW_�50x���$���<z�����±�k�C�}���f�oKBY�kX  .�ٶY<;�5�H��-!�^]=�`����x>��t�����/n&6��RV]]��ك?2F�o3�G�6�>#�VNNg�6^��&��#5p��&�~v� �>���?i�ʽw.��	�慄����:I��������@*�6�f흙�T�üm$��V��BR"{����6�&�B������4�b�萎�]$뱄sp8�뺟c�����y��<�s_���]��}������/Z�}�`$�8Ӌ�b�n8HZ���x��jV�ZB�B�$f����&Nv¡/2V��I&jn�p`P��l�V��c�(i��}�:tI�u�xAa�j�%ըY@�'V|~���a~X�d�ɿ�)��5���r��Iv�>��e˖(�m����c��}'0��n�A��yN��������ψ-��o�o�u�=��ْm�����8��>���5id�ΤC�{����K�'R�����h��X�V�3ˆƶ�S��~,a;*����{(�u�U���4�����Py8ef���nVz������==����?�8 _0���9i5��S���'&&>�3���nrWi��_���K�6��M�v9u[�nK���8�:;�0�g,�R��R��յ}��b�rM���;�-�לhѺ���z�ef���J6��Xl���fy�'�666G����#T��� ��&�������g���|6{�h�~M��;����R�w��B�4Z�@  >w�,��#	Uź�I�vj�5�y�z5<<��q����:S3�0��f���^P+�=�� �t'������AU���J�1�&��r,��*i��vv���iT��@�2��g�����vc&��w��3�T6���Ny2T>66Fw�R+�������EQ�-��ߎ�`WФ��!�K]]����Gj'�+{�˃؊����X۷oI��"��&VV��c�,��،����{f��Lm�]����R��S%�m�:456^����X�h]N��o5-*)n�25ՆB�D��v�\ڑ\o�O�D��ge�}���-��0'ҿ��N�B��M2�����;��} ���Wow ʄ.�e�am��k�8.Jm��l����u3�OQ8C�T�3=xv_���������ʌ<�@�/c��nx���(�]|r�����f�F��Ò�[6�0�̨��X�[h(z
>�V<+��p���3�l+%�y����g���ؑ��ST#v
���~۝1�ma-�A �9,({55�5i��.���5��?���a��
;��8ɚm߄?�(~����f��m]+����ג�&Fo��0ε/�{�uH��YyV��?��Ηa���7���Y��2��mtrr"
ǹ��iA�ܻ=~�s�Y+_��Q��㣘����['�p�@�]�wFY�&�9G� Q��ۉlH��n�dԍ(8��j�ؾ@Ȭ ��9U-]�^���h&)������S��ףYYX�OMM���8~7��l�~���Y��U�tOu�����L�x��!�k�[�M�B=9��l|�r�����_�R��Ԥm��7==�ʣ��Ԃ����;v�Αݾ}s���..۩���{��&�t��L��.ᄐ-�7d���Ǐ���\�&���[�BCCw�ݻw\|F��+���+��'F���>}��f�� dK���ZZ�����M�&���X��6�l�KJV��O�(�o���!�ܟ��S����-òb��{7�I������u>������|W�-��f��Op[y�����.,L��3�S����u�ЗPmQ�"<q��x�ν��[k�C{(R:v��t��ȹ�ؖJFE�������<pkE��������'����:��.BqyQo�'�X��x s�j>��u���ѝ�<����z���[C9����iCi����ᾀ�y��~~����ଐ*d������57�bM}��[�̋����'��NsF1���(*� )!)�5�U�P�Oo�el���@䫔�%Q�Gi�쁴E��B�>��ӊ����,���\��v������*))����Ԡg��!/���w�ާ[�^�r��ο?L��)P;!c�u��) %M�7Bо��]�_�|h>��S�y��<t��ϟ#-����[y��l���qډ�W��9V��bNYg��2̱0:�c��u��Q�s"���Xh
Lr�[��JF{�7E(�ǅ�.C��8;�6�A\] S;�� �v�]ٹV��7�v�3�^2V�h�� \�NZ u"6n;[[���:$kYq�(K
� W��*u���9� y�v�k�L��-j���y`���L�Ie���l�,VgM��F�=R�l�W�����i�Y���I���D��꾜�	�R��Tt��)3�� &8�f�'���h%( ?<�"���w$~hl<�v��9�U��?]<g{!��}H7���x�n7y������p��Ǐg@�T�{fA��.�^���)(q@��m�v)(�T��dL�u��1���Pzt���f�.*����=�K���] �&+����]k����޳g9���C��|{敶��	d�V�z�x�\e�=i��i�	�8�@7���Жܻ�&A|��Z?}
u�8�F����'��p>yAW�u7>>���$�[������~:8�����F��?����:X|@.��V�� ���>��j=,䊎} ��ay2릎�+��&�����Al�@�C�^i>~�x W�wU�r11������ؕ@~������P�ՇaD��0�p˅��ë��mV�UVB��o�lĉ�C�Tfϟ��8�mq������d�ȏy� ?<R�Y���F½{!�FG��������O5��SQq�*@p._0��88<�]nL��g�^��m<g蔯ع�}<��C�%�}�z�H�cU�O����v��HM�9O���q"�Dݱy̶���5��k��$({N��P�r�����\����ળ�����)+(W�#"#����4T"y͍N
M���(��W�]iS��k�o��������SM�1\�7�*���7O��O��a��Z��%�/���w�����.x�e��u�{��'졲 ����!��MUH2�J�ee{�{"B����wO�}BDB����䷝�=�q2��K@u�� -u��$)��3@< �s��?���)(��N*lĖ0��UhM�oR��'��IY����<���-C��޾�3���]"�����jh0"1��S�$�������+��u�[�����A��H�%I� ��/���Ќ�d��e)���/��+�Ml����#��(���B̢��5\�Z;s1nu �����������_kcc#4��(�2J(��
lQB��sM��B������Wp��I�]�A3�����is��'�k��C��4�|R�.��)���/_>���d��)�</��|A^�2�����*�+Q�vΥ-�\w~�'�[=p�g�sg�p�1ߞ�XұDMN�X1������ˤ|��P�����w�o�?���͒�[�
���j��]�D������B�=��7��[殺���P���?��o�K�|'!A&M�0�����>�9 ���s�)5�칧����W
�4h��A�zgGGi###���Y^�V���'Z~�A�R�w�=�ԥбu�� '�)ħ��Un���a~�֭d_��|S��^�9���C���Xjoo�fL}�_-!���.��O�*��]b��f`` �}0���+CjU���ҿ�f��nhI�{�r���K=��8YvN.���u��b����P����k�Q�TpU?��[�{���e�r����\�<�;��qTpg�	5xx��/�d	�����w �&&&px���y�C��$1`l�&\�ȉϮ�����nSH?RkKK��opŻ�]x�jk-�v����'�-�U��"�Jq����ɵ��~��]�eoȼ�-<9�c����P$pK�����PڡE��4gh�~c[ܵb��h��K�n>��������Ez�ڵ��g����[Ma)WU�4� �K]�Xߌ���C:Z�Aq���s	�o0�@���06���?}ؤT3L��o���+ZZne��v�
���FO7��Y��~��N%ԃ���y�j����q.�{�66t�>�^���mm;H��P�i���w� �]\W2��c�D�?���Ķ��E��C�ԃ�_�p-��ݽ��ҡʣ�Rf ʾB`xx��3e��frҷ"���gggg���y�����x&�խ������A���7}��Y���T�Ì95P�F��UQ�1ϗ��G��X�jUگ���������6����8��#��AT�?]S.+(+[\DJ���s�<�f��9x�ch2��O�/�gA��_f��qؤ�o]Od�AQ8�.̀"�*�i�I���*��
���LIU�SΝ`[�*@�Wc����ar&K�@P�1�>|8�����6��3�Fr
�ъ��}I���N�;�������㎊�5�s��Z~@e۳���K>�ؕ �Ѯ*�1?(O�)�b�B���r�Q�[{yɃa�����\-j-{}�F89wi�24���\.��;a{��`:�(�G�5Y���u��d�DF3ù�Om���ۄ�5�ɉ���:���@>��wt�'W�}�
�]`�˗/wd����]h[;�{aeݔ��\�g ]	�7����OL�(�/1�b�����4n��0UW�~b�����m�i��jrR	F�r��b���H|��a��ڙ`_ʇ��@��� D�YKHJ�*��5��슄Qw��[��d)�n���_/U��&�Ru%�K.�@���p&�5p���*�w9�@xd(�h�4�)��� $�#�}�W�.Ⱥ������mi��-IձM�m��Ȼ�$]]w e��X�PA̐"E�%#����v:'dfr�.��Ɩ� ��J�ob�� �Ҹ�q����(���LN�mk����_@���N�x�	�v�O��������>�J\Y򡇂9-���{�؀�Y>����#�����JY���t�8��Ą��}�p��m`bZOI�0Q��������=$���Y����۴�j{�^�.W�*\��AU�����4��ax����1|r�Ņ;�������MV�ώ� ������<;��d��� �E'����ӧ��=9�����.y[笠��
���Nô�{W�o��t2�	6����ND�S:ݒ� ��:���t�һ~����瞞�&3ї������^d@K(���F0� �<�m�j(���<�L�[���n�5#�1"�mK��u��^�����;r̝�֎Bp_@����秱 ����%""�K��3_�-�ժ� �}L�Н��[�:���3��UubG���~ZXx�t����
Z��nL�Jd#��!|q�To�z�8<鉌�f���R���>�(kTn\��m�1~n�;����e���wC�K
��
���\	�`v2\;mt���ӚA�V�O���������DuL����.U�{O��!��%$b���"���ܳ�ϟ?qL���p�V>?�@�_m(�̱ml#c�O�6�Ӏ����!�i(��;����Y,Ǚ�"!W1O9������3�ROs *��66���x�>d�,YEE�,|R���X���,q?DzI%����'>�Uu�$��s�������쟮j��d���P�!�Gvיִ�	,h� �@%AmR��6w`K%q*g�����k����4�3d����EOk� 2d� ��Y~Z��,�Ť.���bZ#!	��ӈy�l�J����4V�'�1��O��z�}��o$�J��#�����h1�,c+��)X�3����R�&a :Ys�/�pe�Ț�?��0��y{��-�����砦�Z�$A���4�c�ɡ3�xC#�]0�!_������ �4�2�i�e��N���U���9���j!� ��F!����!��>����Q2��|3L]���'@jڒ�� Oo�V>:35��_b��EAi�D���)�P���x+�W�Z�z<�v+=�چ�=�nBC����3�J"ԧ���3_�+;�H��wvn�w�m4�L�
f��� ��?���ѡ����ں=[���)l����^�v�H��4��,����95hB�9j{��" �TXI+[@�W��~�6�@��`�i�喰��ɦ"�	�wA�l�$R���ԟM�IU�*e��vZERJ�}g�z���w�b����9�o��ï�#���$p �d �
{��!M,��8Z�.p��=�����8(Z�E�~��{D戄L<kS���{�c��r���pi�]?�ɬ*nV����~$�}! S���TO��fPh˼ǝ�	��f�]O���i.}Z��0aU�Bs����k{��hU����;! L�<ht~UWg@]HEx!��8�b��FB�qR���i"�ʄ^]λ���CXBңlM��*&�!	s}	���Ɍ5b�_���	��xԊA�B�Ī���h'���*���;�,,�O��Y��f'�r�3N�g�^��O��/����ȭt� ��z��V��m��BWo������7��s�]�"�Un��_4���ׯk������̔���$����߆#���hM�Ђl�S�{��a)�Pѻ�~W����7{3k�hO�4��M~��A7��jTand�E��" �	:�l������p�G�h�㸋|�ր�߭���뙙��r���pÛ�ܓ����u�m���B0�dښ��t�0�\�����d��q��ʵ���x�S	�%}�\����e8��Fk�=UC>�,���U_�O#o��������b�ƍH]M䘷��	�fL���n:r��
q|�8_��P���*��Ʉ�$>�Y���Vr�[;r����(ܰm(-���¯<L��ʎ���E�]#Nd�y���6&��e��ŀ�?AM�f�/_��Q�)�]]���$N��A|�E""�޳���OG��ʷ�OzJ��fn�rhȵ9l0�X�f7t�1{{ϱi�}�]Ǩ+eePN9^�wj �d`q�b=y2�q5���3��a2Q,��ب�q,\���c!�o)�s���օm3ιw��v����,�����v8I�!���#��]���/��Z�<(�p�������)Q"2QxzH��8a$P�5W�E�&(����Js��k�&�ʹ��^��	��޽K�K�@:Q�@�eEǜqsۉ�=Zۧ�O�8�>�f��B�
!W�;��~���������t���L�K!j��kntm-;�xţ��K�^������!��ρ���eU��lz��B�nI߹�#F�.�#���ߗZF���E>�m�N� ro����ݛ�(:Na�fg2�w��f��;2��yʨ�9Z%"99����%M-��8���J����8��oX�pa�caS�=e�C�v �Z1�pP�T�&H��π���ϨMi��W���s@��c+�R"@�@�r	PPRZ�Z	{�8�/�]tf&����EWg���l'�ߤ�X�r6���NkL��O��oo�%���� ķ��s��S���^��i�v����|�����8�5�=���T'�����Uu�)::����l�X�
��]��e����嗀y���AZ��h��a���<��`Hdeq��=ggO(Օ�p�͙3�*[	*�jjk�!q�%[�V���Lyɇ|�Ɏw&7۬[����)@AEe�|tFom���{V�Z������>�����MćJNǝ�Q8�r���}�$j��n�z9�����m�Ǭ��+3+v}��_�3׸�U��j�s,j�"�"�C���0!��v������*+�X�`)ǋP� �4��7t6��Ђr��e�T��o���X�	�4a��=	p}�Z�57�:�R��H��8|�$T��SSSw)*;^� �����j�g��8"�M~�SRR:��k�R�$5<��#��5s�w|�����ޥ)�3�\	�g7�b����d�>/*@Sg�#Sm��S�i��8]8�70��Z�N쎗�=	�����8��x8F��"U+�,n����� Q��[	4���G�p�ٍ������M{���#u2�)ː�r�#v�����!ǎ��<���B�s����4�X�JY�%9��
v�l3۪�E�_ ���Z��	�uT���kϱ(_	�pO��,�c�.�*��4ྜ��$����P�,�� �Q��p�̅[ 9�`�����+� �]{��x#��	.����U:�F\<Y \��X��=��$����`���;⻁)"OT:����S��H!qj-���|Z����^�V�����遗��Rě��Y��o����9�g��\���EQ��k��$%�*kB��j�,�fL0�d,�a쁘�knl���lNtqv~�](BVR:E�8�yy~���{ÿ�����FqߟA)[�ؙx�F6�ő'KYJ������[�4�ݻ4���ň!��Q��P�׀Q_�h(u���k��9����n�sju%���������߹s5C?��T���w9;�b�2vO�币\5�"����'�{�4�q�_T���j��Ʌ����<xW���@�27�!ܰ�2���fj�՗/_�z�~=6G��wt����!����1��7{��#
T�i���c
e��t����"��HE+�MT]��BZYӼ�{{�].���Bu���N���$Q|��Wu��*�NUf�"�x��U�ȍ��{Q�7f�+�������5'�1�ٞt��"���A�)z��>�!ssz`� .u��%XOP�Y���z���rV�������߉F�}'��}[��Wc����#Qy���7��s۰xѢ����[yEv^{���E���I+�znn?��wab����WZf�:�*qK�G\�F��5�}��wAC;��-Z��3<����R��kr�6X5&��\K�l��G��GFܨr�@E�.=#���.}p�.55q$Q��@�y*H_��ĕ��]��d��nMMMA����g�����"l;;�N�5�i%9Drv�,�zP����Pb�A��2�1�J�(GjF����.�S���	�6�p���u�7��N���T���4�j�b���FQ��o/^īh�͘�"��[E�@��m�k�Y��~����X�h��W
��8������Qltܒ�3��>���-Q���t��h�F�ZPY֔�n��	[�b�D����ڎ���Hq�~�.
DP���֐�ҥp�ƞ='�o���!<�o�eq���̕H���q����{��B:N���c�&��mj�	�Ŵ��I��]��}��]�Ꚑv%3Qh�9j�D��t�O\8�%IEsS%28}���k)�p�~M�T2�r�G�Jx���,�یՉ*ӑ}oWj�Ml�!rr���zAb����x�x�;4�C�A8�9RQ�7Q�Bn2o�L}���9c���ca��O49����mC]2ؘ�M���m'��t�C:���G!�\N3T�իSSS%>Ö��&1�	j�I��\��gPt���*��F $�GU�=��Vq:_��Ã��:��m��x��t�Gƪy����_����q�im7��Ӻ�J�o�k��|{f���d���ݻ}�
H�4��(�#�}|�� hi��0/�U%i@���������])� �����f����>�]$&��*���j�7
���AK�B�K}=����gFP.�"�;��f�T����f��WVV٣�E�7��k�.���6Ȝ�é��K�8E_���s��J�䁒�s/"�N~�K]?hݦcK����p��9?�%?�߿62B�D��?}�
���y��P�AD�⡇�-��n'�ɓQ.h	�]��
�m�J���6im�o�ݚW��^���㟗ѳ_�0#������A��s�o���̞��>�5t�w�ܑ�@�12u'.�ӡ����p"�d����DBY>l_:���-̷�#n�y�;Ed��l�sJ���|�v^* p�RP��(S��9�c�ri�#�4����5��x^�£JԒ`O��VT�t����l�F��V�G@è����j�i	��������$YP :O���]��bRL���7lW�e�Z#fstH��*n�CzJ��u�&��3��7�𗊦"Ui���)H ��|{ �zV`�8�*��4��xw�
��gLŋK:��߼�����-X�ҿ4Q�..6�&��г�����vws��:��mIT�[v$j:KԦk�>C/��3�#�T����QAȡ0���X����'�_UU)���f5��3�%�3{����H��"�fRd���f�;	�����������}@�귔ym�{߸zu�ڵ�!zZ�����/�s�՝Ri8��uɒ%��xqhf���-�6�VM]V�z��MGp��f������Ȕ����|*�����g����+：�	�P2L�3+ܙ����dfŪ�/�T�`���\鬔��?!PxfZԦ��?"����K
��qp��q"5�!,�L5U�����66:(�ɉ�Z1"���9�EDp�a���~+"c/oy��hNy�1�6���;i�ˁHhN�����O�d�,ߔ[0��<��� �ɿ�>����A����l�BQ��������Dko�����CBu<&;إ�aɓk�v@[٥�n�}���)����c�%]�J#��Z�ۚ8�hZ�����O
�è�~;;L��`���B�C�pjQ�;jMq#>))r����2!LM���.�<��]8N[���5�F
E��!e���*|�.UU|*z�2}��<�{��J�'{Ī9����79��B�Ju�k��chGmB�l��Z����(����]k�l CaE��)>.�?+Û�-!�o�Z!ur�5y�3CЫ�5��H������
E$�n����g�k��Ar7	R�U���h7�'�R33������h":����rMJ�=���9ei��R���p(�z5H�U	z�Mėr [�KC�F��n��(�}��ɓ�.��u���Y�TB�!��	���~`F�
:�f��i�WD���|> �օy^��K�.�X�i(Y.��$WQ�5��F oh���*2�tHi3O��65��/��%����{�?~�Hɉk�:�>�q�m�H���1U���z�\�u���� v�&�M�FI��X��u� g���5h���5��q�9~���Sb}�����B}CH��[�d��/�q��&U+�@�p��gIj�)\���:��)V��*�ѱER�"N�E�5~���d�_���{�Se�����K]����=�uߑ��'�v�-9�ä�N�c�Z�۷�����-�� ��}�sM��H�󑓱�a�D	IL��Lq;���PBth�+�S��s'>>�U;n�u��t��3�����h{��MЎ_:���Dʽ9�V�-X'V˨a-���+��k4h���c�Q��	�.�<��s��q"6�D��S��."Nq�%El�MG��c���K�����Bh��Y�q�UҥF�8x�ࢨ�`��]��6	��<߈駨ج�A$�Pх� �w>�3'�?�%]�BBǸ�݋�����/G�����(����v3�5@]���D��G��G2a4�56����
��񧥥|��q���з�
-k�c�MNN�/ŀ�Ƈ�@~h�n'�����.�X�Z���]2,��z�Ğ����\��#Q(�dddn�>�&8#u^�ג���?�J�����1�T]_���w��s�O���� �7oR6�b�����^'�:��N�Z��#�P���LЭ�ˬ���.�.M�n�o�d����b��EkW��n�����a7oB�����.,#Mu�08���8Fpd�C,k~όq"���5@�T�Q���Ή���knlhh�>}�����$�(h溺��ˣ��6\�2��4u�l���6��h�o��%wsA��&�N�f�s	��PK���V'2�̈ ����.�G�)v+ձ�\%�r�&p�8����Sff'�����ֻ��5���3����p�����C��J�{�q���֖�sr�!��	�T"K��(qN!Hve�i���0V�����ܾ����G'�����)a�o�Z����G������&�T⿨�����~�������U`	��U.�8j=a׮�x-c^L��Ν?��ݻ��혣�xn����b5v�����X������wD����'ף-H+�o�Ɨ!�3(x$�Y�.����6���f�����R���R�;����CC����Ū�S牐��{�������sr^e�Ƞ�|f5փ�j��������fq�[��R��ǖ�gMґ�ܾ��?4�StŷX�Cm\�g�|������	�|���Th���}vz""_��&9����aj�)R���b<��>C?�x_n�j�s�b�24 l�0 �T�L�Ω�w�T@�'�G^�+O���-���^����kD��{#�����>�G�@�-�t��X88����~��5B�q��_�6���kB���>|� ���@VW��I�^ F)�j��HJh$�y�U�JR\:��a����B����5N_l���J5R3Հ
�O������?�����2Nx?r�������(ť��t߀�N,}'��p�xg��VXJ��=���Q��~�dv���lE�QE�TG\�]�@�&E<�E�֯_o�J�[;Z-�xj�9�RZ�7ć������G�l1�z�nS��7�j,^��H��a�z=|�.�tH�:��D\��e�޺uKU�e����M���#Y�����+�.�gB͘�iv�Ӝ[�&gM�3`<��[[[I	y�K��k,��3�_���'�j�u���Z[-?��:�M��|݋���+4u��j?"d��S��	m�.Lp#�u	�˸��}jj*τ%��]T���˺u��恎C��k�*��^N���S��N�ݱ�\�i6WxѲ�GDQHR�	n�|�D@;�`:��|�c!X��V8wy��O~� �]�o�ћ�i��U�����[C!�͔P�n�kǋW�4!B�bi�x��̤���=����nʭ���6+>A���&1/��9��EB0��;pI�{�r��}A�P�e$�Ɂs�f8}%<����O���i��+�/Bb-d�v��W91��9�����!P��
�F�k��l<������"!	]-.>�ok������'?��j/#I�>xff�xF�[�.�DC:��S���t(.��Ҳ���+Ҭ+��{�#��0q�bݿ�wW�LU2�u�ĉс\��y«���E� .�t�F�X�&�fdfZ��L~�]��KA�Ҙ ��klFi��0���&��b�`�ڜ;����>0��f���!||�CO�:��@�[V������o�i�43df$�<�E%2;;'���㩄Tp��W̦#3�<���qF]H�6Z�{V�1���!s�s ��#Q���R�_�L��e�\����(� �(20�8)(+qr�p2�����QF��ܻ^�/��2�4�vp�J�4T�� ��}y�X8I��0
��������E��Һ:::.!�V5m���'����Em��j�ά���B"�ԺS�j@QUf�	�s[e Y!$d�Pږ|�߆:�
�3�<�1�5��BVy��u囲k��� �#fꚔ�p�*d��V�D�к���cۻ$�9��M��sP����q��#��[ը�L��1(���m�S�J��&)�Vk��L:���Z�=�x��27��i���		ھ������H��\��ƾr�J�95 r������J3�>45]7�bq�xYV������ގ�ڕ*Y^`�|"C�%v�ŋ��aЌ/?�I��,���(�K�koV7�t�fq����K�'z1N^��_�K�T�)�?�(��}N0�ZLl��d|�#T"��ŋ#��4cl���D%&�swB.q�F텲p�
0����(OP���״��m�g��c�������j�T�[��w�_��N�$�
xZ^��u���V�Nb���!]}}���QA�,��9-h�F�%�`�Bf�$��  q�S��7{��<����e.�לhUz~s�Tw,�RU��JHU��}6��l&�_ ��ԩSWKKK�R�;�;'<3Z�����Sl�� ��vT �D4x�6?&��2޵sgm��V(��==�O���C�|��C#��g�eC����ތGH����9A��Uf� �c!p�-n,Y��W��2��V�������
 q�~3�z߽;�F�~	�L����q�rn�j�鬉�wB�kK�R���2������(�l��_T�*?��C.ke�5���$��ZZ ���p����1u������^uj�R��Z{��tv��L�)����M��<�'S�|�#4��7C0�dی����8Q�W�v,8�����ƍ�b��p�zzb�r)�io�Pl��
݊�c�C���I������>�R)h��!�� �����T���c4���DՁG/�}iE�S��Ӎ�\�_AV�f�L���qsۉ��l�����$̰�0�%��I��k�UEZ�!�+�2hm%@�}�;�[��oܹ Ҥw��cv�={6oh{���Z"2�^r���@	:::d)/5������C�A����
������
�(C�mp�yfz w׾}M�Uh]9���~�	d�q
c�~�^�M8cS�7fg�WA���&�(�����z'�B���ljr�s��ZZ�	D�ײ!����7���<<�d�`<�-�.�~#�t�#���p8��sA�`��k��<b�?�1Հ>���!	]EX����"U��a&�V-�T�pǕ�_inq5����ߓ����Ɋ�n�T�F�ڵ��n�Ƥ�\�q���n�,hQSU�cz��-m`"ll�*��}
�3�v@A�^��v/��>�d�d��G�E�{�����LN�%�����(��~qI�b�C"�N@(�/�d�������jM��)�z�.��ڬγ��%˾�jxy�F����C�7��ǥ�����V$>j��$O�Xy�rlOg�����Ws�s��J��{b�9������5Į�F��v�D��Dل�KL� h`|�3e�ЭsVH<'����Av�"	�j����;^��Ƶ�a�	|�	G~~��=�0ҟ?Y�,�.7����Xd;��MCN�K²�2�/��n�A����3�s_��J��J8��Ͼ�3��gB��u6�S�RL���ԙcW'ck��m���Y�d�k���� ���B��Y�f�R��99� 8�U˄6�n�$sy����X��7q���FZ�-��A�Q`�"܋�Rt��n�x������@��M��D�P�b���%K����� H�5A��ɪ��Y�|)ܞ♅yG-ɵ�l�'� �_���3*��3q�i~��nE�Z����%�xd	�[� O��-�Į�����U畗�u�����Z�Bk��r@w�7n��n�읗쑨;��5:�������f��6] �7˘�N������Υ �L%�M]B�v|�������BSUn�p&�ckk8�O�D�q�:��퉻�*ב��2�M����:>���
7���"����7�"�?CB
�mM�]\PL&%EA'\= ����FҡJ-���h�׌�:kW��mW�nI�X憸q9+�2�j�qI���,��d�gB�0QWiE��_��� �6�A�ٽ�hv.�2��j</oT��9�2���Ep�o�1�匰�	���О,���TE�#�LB)GN��������M$�BO셸�P�6�x�1mI�Ԟ8����)�ە��j�����)3��S�Rd�Q��p�3��Q��W8��iǯ�-����&U��8ea��-(��ړ�Í��׬�2Sr���5�+��y�H�L�܈N/]#��f���?�Rջ��L�)(���ڀ�q%�(�c����<ɤv#���t��|(��A)�R�$��T�F���ف�5�6�~c8�"�� �$��u�4��u
��'\�����N�7$�y�������E�)W&�py
�Q#�V"�U�4N䎿!I�Y�����E���d� |����xr^H4��w�5�Z2!����u��i8��<��ׅ�o��F�����'��\=r��%!�Q x��M�pG9�7�W��Ȱ̭�H�b�~���^P�-/�b�ƍ��s��x��wB�#ʶ
	���@�:�N���ϡ���ȴ�������m�ۄ�,k�X�?��F���N��<wF:aNkn"&5ۧ�m�Kh�Ϟ}����ˊ�Q��z[���h4Y�!1�Z�B�ş������o���,E��E)e���.Њp<�z�9�O�	��60�"鮉=p'�)�`@M��Z$��1�@�wB�q����߄=p���9I�<jg��X��z _[��s�O���x�h�dh����ʃ��!YYA-�r����9�+��X������
ߧU�4� 111��{A(1B���c�0B�3=�Us����A%�Rhx�b�L��.A_���R>����Xx8�SjN<q�`8�W�}��Bכ1<+�?���>�hH��՞�{�O��7m�������&&�W��(�oO�g�����f��c�<�U����fѫW��s�*F��<����1m���N���������C�U?~gQ�k�ѭ�孠�C�m�"�����*Jp�a��[��7�ڰ�g(J����M�%��V�kN�G~�����S�L�y'��lM�h���I�t������.b�}i���h�F��T���絽����G�|�hAǽ��/A_�8��ʖ-[D�^��2e}��Ny�ʰ���!��???f~�����t��~��2r ��1����Fg#�,�Xgu�V3WZ�pm�$\�w5e����i�A�F������o�4��f��	xe��)��A�L��(t�2O������{�1�%���eH)b�e��\����N�ŋ_�^p�kw=��K_��pN���Cp�eXX؁ȱ���z�V�L�̚ǜ�����H���57%�>;�����3zV���E����GF�����.���3�6�ˁ�����H�_�Z_X��(R+˘I��i|Q���a81��B����r�w����}<g�Q��e��{��}9��љ|�0H��U]"ɇ-��1��uk���)��d_�;��׽�C�>���⪏��37�jErU�I��]����67p?~<3�-f���ha�|%h-��gJ���V�J�,P���+
l+M_}����-�m:*�l��#�XAk��l�<T�zµyLdWz�r���
x$몒V��A�6�[�����gV������q'��-P���	�K�� �ٓJ��Y0�+m��L+�~M�������KbO|i����2vqi����'n;+]�ƳVY&������{��r��Kǥ�������[R1?e�G�}�����ܜE��?���d˂�P\j3�P3<�'/�4g[;/��Sz��x�!��'�`���3��C,�y|u��WNY�����ȭc����������6+�hȾ_�'?��?�P��3����2���ZN�W��
�D�@���}������V_I��3 �C��> �`aԙ�k׭;!����:���K�}�&��{������T���4E�E�	��*�[��ݺ'��m[ن;b}*%Z!۲��_���lZV7�U�⿵{���ѹ��K
���1/�#_qt�=��i�������S�K|�z$S�}{�O7g��6T��gܪ4��,-������_��}����eDF��v�G)B/Q%���֢�ۅ�!ML#� h�;VZ��ip텠 	f���5�c*wӏƍ,E�|�vZ�t��6������n��ILZ_�CZ}�}���e���E)�8 	�������^Tu�m��V���~VV@ℊ~��F���m|��@Gq���X� bҵ�d�����o���ɋE�i�\��d����^��)��߀j���2⒒�` j�*VU�{��x��e=�G7�z�sQc���;զ�A�e_T�S�$J@�>��ߴi�s�7L�)�Y!���_����z�x�JNWWO��ae�c�(����Q͹Q��d���a�1h����|hy2:x'�-�K'g��%�uRz�s�>��+�����c���)�6�šϑU���KB����CT�]�ee��â�AU��Bշ�tO �AL��y�ZU���
�8�v#*�X"5�/�	��lVCC�9�ut������'>�{��9`�cR��ѽ�oa���B����V���ϣj������ ��Bc�Q�H���,�9�Ue>�%�Ӝ=��q5� �t�X�0�C8��7�����Omz�ۜ�2��5�d7/�a��/���XYl�#P%2c����b����P:O&�!��b�Sqf��T	r|�Q}CCC�ݥ���-I/ܰt20Y����m��(���H1곹�������GfŮ}\N�XqMk��xBR%eee=S���6{��g�c֩[�	��lᘊ����#�������cd�����%�5{����5�͚��Y�l��
��Ȫ	�
x.S�Ͷ掎���9WW=$�9���B�h��<��!���!N������H�U��-������h���ր�D(eF��?�\2?�%��Ӟ�����j-�AZD]�r�4�>'����b�'�d�f�ɓ���X��_�8)��XWTT�ɯm�������z�}j�М���:���¥߄����t��珏��c�x,�/�1�9V|�m5 �)O��*4սr�"�5W�
�
9�������WN��wԷ«/��58������[ /х���׿���*9E�pߩ�]��c�����O��ޘ���~B����De~����S ����9������YOy�L##O�HJ���H��g��Y�,qnn k`Ph���..$�I��XƌF��U�0�<�G�8A�E&�z.�c��1����p��c�9{tO�ٳ���N�}�
r�{�����r�fP����~i�ˢ������~|�67�"Lc��7o�$���]�]o!�6"xϝ�0nsP`{A����P���W�1A���GG�~`gg7��0�Я"ө�����5;'��M���+{9;�#��VO�ܧѧ4��?p�n~��%ɸ�  �]݉;���l�>��\�U;̏)Ļ�s�⺔�jk��g�s�|VE@�����غT-� ��wo����c|����+�q:m��� ����Qq�!��X|͛U��R�8���rx.��5�J��~}do��y�"�c#h�{{=4���P� k7��\��4�����g���$�X�ӷ����q)"�m��C�Q�v��#9t�{ 8$$��IA���ƛ]�ܔC5Qy��JX���o�ud��h*t2��X� ��鯥ش��'	�%�ss��xA 5�����-���ܛ9z�;������c".~~��EdF$u'�_�#w�Ki�{�o@���'����kM�~���t���é)� >����V�f�1	�/��I��ҩ��g^�U�y?6�O���u�I�)�O?��
�?ܽ�f�E�Ϋ���
K���C��G���L--!I"�,z~��)T�L���:�;^{�Z03��6T����[��d�}�����p���i)�3�f���䕕��3�%���@7�u�V�"U*
��/�?:��i�ZJ�������0��t�2;`��i*TMb{u��/�ʔ�5�?�U���Te9@�UE��ҁ^^^�jN1�
T�mmm�H�P�-���0���{Z˼t~��'�r��c`�N�81=T>\PQQ�3�Y�֭wP�Ba{����a�,d�caS�~��7�T��g�]}�\ܾ�_�a��`c� 
����e�Sy


��C�8+�1ؕ��9A�\=4�f��n�Y��bv匜W��%c1���H3X�Rs��㍣�`��j��}��V����;���w��2����V���V:lN�%Q��RQ���19��Oٲ�!$!4&�!��(E���`0���<����P����������_�l�������������� ��tu	��M�j9=9=33���F��?է(2*9�C�F� �A	C���[5.��Θ��vd��?_f�}���f
����*�U^ً|w��}�w��'e���*��4����weҎVz�8xTI�y�zd�9Pe�AUƹOh�R^z�I?�3�-���4�� _�ŗb�?��xb�
q*jƠ�41���UWGq�ψ՚z�'00�TJ!̆��1c�Ur�A�J$7k�7�«�C��xj��U�'��Q�6��-�toA(�����Ը^%��I)�Y_OO2Հw5g2�Vr�'�*�ׯ�C����j���m�74ըI��.�3�T�Ȍt�X�I4�[n�H��_}h���h���
vZΝ2�������+���m>~~t�&�úk���uq{9`�Y{��C�������A<�mm�=а $�F���Ǐi.��!Q���������<
��.�<!���aRS�������L��R`�a�8nա�lY!��(�m����-Q���Q�U��BX
�Z��%�@���RZE��R�՛Y�_��Ga2�ȥ��rroBNp��w��,(���y�	�B��Z�D��>�?��I
�(���u[*H��}�US��]�������*�GJ,��N�<8�Z�z��2�����fK��|3����Ej�FY҇�G�G	��	d`���R�b��y�!�[�1�x�NUj�Z��y�'���9q�2�UP ��H�*4x|��άf���8@|�Ai�Q�l�i]�؂�f)��ԃf]I�xz>�;y}��Ǒ-kx�����6N��Of2��f�kv��d�k�A��r Q��Z�������B��zȂ�Ѓ�7�6���
�"�Zi.�e������Ku��K�.�c�X�h[K`���ONNV�d� � G�f�Չ^�<���`���p��� ��䙠��s�/���e���H� R�h����%$�0�N�����b@a�W� 8t��v��s��(�����@U�L�����8 �U��C_ݙzR-�x!�2J+Xʳ�!�'ԽE�|#,�)��Z ����~!>)!�2iot-ѧ"�e'۬)m����0Z0['2� ��]���j7k�KQ���j���ՏQ��,��;'TBJ�E5\H�`K:nd�_J�U	��}�Ŷ$PL����(�(j��%4�'�v ���(��s�k���P��?&A :C%���>}Zߖ\j����\y�2�Zmmm3�Y�FY�N�C2�TaSס�C� n>%�5����*p]of��������n�V�:��ф�ڪ�Z�¡� �<xpx�>��/�P�-����wC't�h�Bm��J,�R+q�$�
��Lp�({��-a��enn��&2����G��گD�_���ylU����t ��@��sh�������<�������bb�5Q��J��}uq����s��N�}����3�"Б�ѧ�:Zeh¥��6!�}�H韯e ��P ��<��R~˪��i_�F<�ؤ�~��i������2jc��TZ�-�������P��~��L����a��O�8 5�S�F�ŝvS%UU�`֠ܬ: f��N�R���d�]�B�����N̨�h��׍��6�Y5��x'Zw�X� {����e��o�n ��}��]�!X�s1쭲��/c�/�+(E�:��o���u:�6��t���4��&��3
E�x�)$���D强��k?[YE� ���@kL͍�&���4ܵ�݅����D,�WPȆ.A�B��c����F��F:�Ç���H�,��L@4�9�zS���C>�Gj����[���.��{���7o�xg��m:	J����jU��X��P:��{�O����s�?�EB�@���k��}fFZ���*
����A� ~b?Y�ȇr�M���Z�AYu����Yn۶Q� �,4̤6��9C����W�`��U-����{�S��+���r<�D�rz~0a1P�CY3f�م�H뻄k����9����)�����˒|�6�d6=7�=�vXkσ��gV��sj"���^�j�{~;+��5h�V(����D�lNe���J<��1C�%��ܩ�����2��RQ�]�Zv��ս��SuŌ��v[+ެ��L�ooGLS])�l�̞m�s�nDD��'y/<��f�/L�^�����?3ܐ��|��ͤ�w����D.)�w�����X5��nr`��ީ��p�n���ǪJ�KÑ��Y�DL�`���_-9��795���۷7cpW����6�?VI�g��H:**j?��V�%��Ol�y]����h�����"u###�ih�|d���2�����	�1cjH��U�^�sYs]9
�T�C�{��ڵS '���~�V� pn�c8D��k��J��ܳ�"� �nܸ87~P���:0��6��Y���2T64P�l�����`՘���m"�ܞ��&�ƧK�!Ս����/�srJ�	@�;����U����5P:1"���tM��g!�Ŧaˌ���/���el�/ P\��zzH�iq�����1T�ݭ���GF>�XE�������j���PN���V�0���y�NE�2޽�|���if^~�������Ix6#��`������.�a�7����tF�x¿��q���:�%>��t�1@�D#]S�R��b�jhp=��Y�q�RՇ@� ����8��<T8�|@`4X��k\^yy����3�P'����g������r�-����fb��J��:���g�G���0O�@��͛��.��bOOd<����Xg=����'�w��:8)\y��пM�B�;4:M$�ڴ���vp�$;c���]]}��x'��|��!J�#ǃ>!t��҂�����=8-�d�B����+ ]ez��>�u���.\�h"S����!�C��9�P!I��m閖��r�s��~Y�u��<�֣f�����	�Pq�|ɜ��/n��V�U�=�yt����b������}4c��C��.�.������ԡ�L��(�2߿+�vCVJ
\���v���Gw��mW�jy`g���Ή��GP��i�[�kxT�U�h3�H!�L��9��J��3��?'���8wz>�z�޽7�2�9��n\)�<�n��S��!sݱs�_�?�_� ��!w``���q�.��T�7��D��[*ξ�	�mu7�>�)�%�{w���H���`�+._L�� ��C�|!g[�'��N2��'y��ݿ����ͭ��>���؃tAX���Ha�0����M)ĉ�����%�}���-m8
aL$"r+IO���-[�0'�::�J�zWP�Z�5k�ق�����Y:rO9�F�@
uDH#j�3�P#bX`ú��=H���ڴ�D��Y���-�Zr���d��/����X�����S�������YK��!��1NHHׅ@+�D��T`���d^)��ƣ�/u���j��ﳜ�y�YU/��B�O���s�r��ٳgU��y[��>�=,sh	vuׅ����2.!�4aAc��r�� U�*���=1Y��'9� a?�{E�y'v��3[[JKKwg}P�Z�'=��s,�i��UK������s.)$�zY~�u�8a�X�n���H~�5e$��f3b��T�j�� 7L�����V�m�<��אg~uź�@YF8�|_��L�����@:������{��kG��f�Y��b�b0%je	k�^��Eꭍ9������P��QŴ�������ڋ�����g����Y�莬�2�(�-ح666���d68AlwMX嘛.1��� ���!�ckk����%�����8?�X���`L��!A��1�~��A���ȷkG�	 /�X.A,j0vR}=�X�,�O�n�۫&)�n�:���ܻ���\]���D"����|�]�8k@��T�����ذJoϠ�*9_R�~�E�;_?�!!�md��	֬}I� �@`�J��/���S�'q�V:��>��R7�b����.NN�7n�P �����܌��IzO胕7���V�!�{%6ԕ��W�=�� mR��pSj��/@�!�_�<
Z� �t�f�*|�0$�R� ��\ɦ��RZFF�����v��ȡt����5 �e����<�H�V$}*����c�b}�,m4mp�z��D�M/��UB���3Y�?���� �������{��*;Ҝ���4�;-llH]X?Li��7a������w3.����I���T3��q��u��*���g"aMI�ǻ�&ءz�,v���?Ӟ�h�����iƹs��f2�K�8��`�� �I�X/�y�r<��З��'i�A���i�^���{Xfa�I<-˸)UՏ��r� n�,��$�Dי�f�`9>V1&E�����%���مN�ȸ���$��/d��������226Ʒ�=����d��쬳��)$d��{_�; ���Xh�D���Ҏ�4�`�-OD��w��b�R�=�h�>�p���'����� 3&&���p�;[~)ZS�ӱ����.q�ϫ�Ӆ�42օ�b�۞����/B��YSs��e����]�<=�8��q��C�����w�ۭ_c��o֯�9>B�>���U����ps����G��.$�xA�ө�oL���U�^lJ�,�`���ަ'�΂ȓ��3��mDl(G*���q�J����R���Q��ʠ4�q��*���h2��^�`s���wW���*�Xl|�}�Aμ���d�����J�fy���3Y%y���Wa�??���a�s�H<T��*�`���މ=�K����K�3H�������q��j{>�+�#��d��С*��J8�:�"J{�[N�Ò94�9; I1����&��BAqh�W��JKWN8�b���eX�ѵ�S�x:� g���;��q����Ȇ���v�ٱu�&�+a��q�Y�T��J�kԁ�BƷoO��}�Ť�R��fł ��C~Ph;��	-F�����7or���t|SG�b�/����"m�5dk��)Dݩ���k�9T�'���cqk�#��*!ZJ��e3t�|@��E��[�=�(��4�T�CMرc��݃�� 2�|�7���E-���T~�/|��R�P��lg��3E�)&:z�3��E�lW����?�IZU>U��AC�?+k_!l�j�����R�'�.�Z>|��#����0�G������dƹ�Ϲ׻g{Br�O�y����
���:P�f��o�'�������]�'��b��\���"�Zݽ�9G��=TS[���C���:[�I,���ܼ	��W���!6k0]�!W�27x�ÁͿ�ִ���N9Ě�ۊ�({'|�ECaH�:�����,$ࣨ�Ekkk	�\�0m������	4�Vk��^_gW�D�(����c�̅q]!�O�z<�x�?���~-;��@@_��2�B0X�5���z����o�9�^\��� d��8������ �E+i���mRx�B�Ň���=7���/��>QlHc|HX���6�l�[&=�L�>C�v�gZ-�P?JnѤ~������dr�UB����n���� G���k+��xv�}T�,,,|�ZWW�����]�ڑ��N��ǟ�8;��s�κՔ����q"o�h�䓳�}������
e: E�BP��i�Xա	�r��~�@퍕����n��<'��#�W�@JJ
}���.��l�Z��H�h��E��v����	v�*믑U?Y�lŪ��㥥��9�
�*n��#B!�EP�wf��ː8�2&�!*A.N��^�1�	z8�K/�Ď�b)(F��b�� ��M�=m��F�yK�j�����-�k� ��N���x\����-;4�C,���[�d��=ˮ���pK�U�5�f��ҕ�̀�G,���.;����'dO^�{b��e�1��Re��!s�6����G��I4����<��LW�����V�=��� B���Xd}�|�Ԑ���;�����{��5����W��߃Q��KKK5	��*��פ�]�l��o>���X\[iW���܄-�������^����s<D1j3�0M�鱏#~���'~��2��^<�d�1�-n��G;B(faaa�A�*�	nS{3��,s/�A�khh���xx�b�W��1�@d�X�E?wt$�Q����1��GV����,���'�������k�m����o~�F��H�\�G����>��O��6��8�ߑ�H�3�}�nD��{�~N��[D�~5/W�Sx�5r)XChg�b�����g(ꉎ�oO��sW,�5��6/0�ӥ�X�0h�ֿУ{�3Bػ�W�2�Gw��[��P�ʟ@�=��V�ZݱL��5k �
 y/!��	�g{u�A�����'Z���ީ=Q�^X����"S33���["���wN ���Zk���E���"�������t@�Wϋ�J݈ׅn�2^�}Z,��W���t�9ͲJ��D��%���������ݻw�U�	�����tuu������
~�~����G�s�����ld_�ku��L}���o���>�g�E����633�6)��\�o�M��E�ʗVZ&l��s�I%���N":�0��"fR{f�O��La�Y_���z��D6o޼�Mz��&�N�����CO8��+����9�����Q��-q9r�)|��ʭ�g?dCqA6o�mnLa�%\V��g�r�^r)xնg�'����$H>����L�ӷ�E�#N �������EF�;����}� >����v��}���w�=��F�D��ps����(����udĘ��]*��x��Z�/�5H�aA�3r�QJ���V��X��{�h8~*�U�jY5c��=.�����<>����T�|G����U���jڋ*(pvs��X�h�����L`���!!V��Qn�QM���g�El�z ��En"���*?�1�{��4��z��D�w'�l�/#��)��R\�C����
�;!�m��yV��I��s�~&j� cdu�@��C��֫j��[<�W�'�>9�rҷ��(�7o��<���<w��	$��2 ����"������J{rrU��_��oA�d�<�r�I��F[[[^N�:T��i'["��"kb������n�Yw���P�`�[�+��&�?�{
/�����j�w��As�wt�+j~%ux�5���y��V����kv=�~w�pb	���4�g�E�똕�R�Ђ�,�~�wYt9���W��DI�TM�TU��p�p�����!<��~�H}��e�w<
�Cd1`)� �,<l��{�� � �x����BV]��0Pom��0!5Ig���ɚ����E�M$��h#S-�]0�o�z�J�h0�z��CD�C)�J�p�U�������PD�P��HF��6ke��@�̺mdg�o��h��fTYc��Ǣj�[/X��1�hWr��U�&�<�z��Z�KHHH���`$O�?�~�u7ci)��/�?V+��}(�cZ�]
hP���OC]�z�ָ1Pmt�a��Har	�6�gѦm�喋���8�ѽ�N�^��o�2���Ntf��h!��
� �/J�P�����Hm��m����j�W^��+�j �j�v�)S1#�y����U�'�ܷ��}[�) ���}�����l��i��DQ�ט���i��]�M��ˊ3�]S�5�Dc��������Onn����9�' �PO�R�V�w�� �o+E]����8�����ё6q�� x ��@|`o�W��i���n�x��<�P�>d�+��HK���̜��3�ޥ�Z������Y�!6�8(�����M�p���(��Nf'?��טzR�FGP��c�<'����S�&���Θ�4Ͱ����n���C6�Ц�QSx:��D��n�'�f��g7�K�K�$G~�N{���jdf���������^���������(m���Z�?�VTO��yE�	D��&�����l�/��%r��-~fU����O ���@Zm��w�&�T2��^8#DH�M0�[*���6��{E^AŃ���sm�:n�U^���������b����t~���C�(�3��?�M����+���%!.^��� �(��_<���O����|8'd1��:��5hb�W/Cֺ��u� ����9�R��;vm�SDj��C=�:T�n�(���A�4:a�Q�<�C���K���zj�"�l���)��y�M�/$�iCK��E�0�D�yB�����(ӷ�!����^8�EKK�(���24�>s߀��dv� �et�ֈ���ef�M:�.8��Hµ�,bN�����ߣɱdK	��P�YYA��u��g\e��JJs|�Q��#i���#�3�t�j���M������!�!����м��Z�M�i��ƹ��Ad[I�ʃ�� ̅�\ɡ��T�w>��h��R4T��ԙs]��X�4�M/+f;!��1�	�\���Ѓ��v,����E���\�֝u���Z���~[��~�*�<r�:��	����Ӆ�����6�-��p�v��`�?{�)�����߾m��%�z�u�w�����O�oX+1ao���H����ȍ��ڪ.�z�7��&c͆*>݌%��痑�/�z������h臦������Mb�!�惛'^�4�D�GT�P����+gS����A�o�$��փ~��l��4_�nUY}t4��H�UM�ު�Ws����&#��G1!��K]읱�(��x�u�f�y3�Kc��v�4����􁹹��uW�v��3����g4����sX����?8�0��~�H��L&�Ҙ�g��)�qZ� (��1�N
����=��,I���(����tx#���ӳ�	Ǿu�*YD �C���-��IYC/�MOK;P���ӿ'�TFN�f������y£��s�W����K��eOx�B��ҟU�Vꌗ����#}&p���]#RSS+g;\hR���	��&�t�cb�/�(>��ǝ:C�z ����Ü���̕{d59>�F_l�����4��B=�y��������|||^���x�E���Β��_�&��s�_/�J=�k�ܮM�1aj�r�7���'v��"�+k]S�����o�3��ծ��JTsI�~ɚ��%��r �0=��5g���^����� e�
I���R�I�'c^��s�)[B����՛�zì��MSJ������W:��9g��aUUՀ��"j������sZ��Tا��0�O���Ŧfff
	[]JiD��Ѹ�՗Q9ŢBB���4a$�Gi����Gw��]���	D�a���O79[��dg\wm�u�8��vO���̇�A��v����W/=p�m�������h~������Yb�X�5��p|����w���N��G9a�}5S��� i��e7<=��}�v�K�|NN��1�ʪ�D��`��3��۵��q8\d-ȣ@\wv&��\9�<���� {�v�L�[��Y���&&vj"�2��������0&&�	Qi�P��tгN�#8+�r��t��gyy�]��c8�|$�ʠ˝�*�ڞ�ե�$�<�� �G���$?tuu�����*���Nyy �!�yyg�H�g6?�ņYk.W`�)�°#{Y�/U��,���7�B�j�7ʊ��SS�R����#�]]��k˗ao9!>��=��DVu�}��2�<���3�&ǿV�Y٠L��f&�u�b��+2�y2|TR����dݭ��:�����~i�K5���RVR�'� �{��-Qa�Y���Y�	��Z<�;�{��0��g�q�~�����,�Aat�`���չ*`%	�9�L�+
��U ���D�T�#P��X��/t�6��V�&.9�\�����Pl>0`_l���j,�L�f�"uФ �ج5:�$�{4��8<�ٸ]�Ѯ%�n՟�p����Z�}"s�=r��������9�Ο��^x�����t�������H�~s��@�ol�(p>�6  G���Ȱ���Y<�D/��d2�<6}�����[��(�oe�`�9ͺ9�uZ8ժRC6?� YȆ�+N~�2�2���l~��i~��|��W���\&���@Y�ϓf�lbe���2�>��6Cs/��,TV����Q�.�ΙO�'Qx
��s����/�;��x�5ZV��fk1 6�E�d0�`"1��Pk�0�� ���)����X��3:xi!�����NO�@�������A��e)�U�N������+�����[ ���JP9?�+I��	G=Yݏd�kznU����������?vK��nx"ܰЏ�K�޿#R䐷��9��^��7_SI��K�V~���Ð��pU7��`]�İ���|Pĝ0�x�N�����&&�q����Se��3�HE�A:���,>5�W'�x��?��i�h_�Pd�������<�Jq;h���~폘�GA�PVV���Q�LN恐��籶9�F�b}�7�>��R����[}e���m{}݆1�*���*GQ\!�q�Hw�HYjwh�5��H�)�[�a�ҵ��u�>;�����\�&���:�#�˃Yo���z�L�>5���s�9�B
��t"�����ow�l�1B&�#ȡ�.w������@g�)+Rn��`��n�K���a"��:TK�S1�)j��x�)�:�Ͼ���c4��I�kUz唬���T�0�!��,.�*SH�-J�6�'���@�候@��ݒ2���WI�761��OL�i�,X��5�⡒?��Y��0��1�ẹ�����H�300�
L~}��9 �t&��h�/�mw-�A�E42s�&�j�$�M�{��J�|ͺ�"Qa\�)�\��"�i~�W�Gps�|��EP������ērR�>l8�x��������)��KƱa�uC
��h��&&H\�"�����ף7����f'�@�_7d������s�R�bBNr�a���-�O���]L������Ǐ�5�3�0u�w�P�n1�>�Z� �@��Q�[�$�ngJ�|K��Yʆ��P1K�x=VV|�۠��<k�֌�Ӊ��8R��  r��v�����hbz�Fg�4�3��[<k#I���[ϵL�:1"��Xу�I��Z:���ųeIN� !h��kgn��6�oO��+#+RR�=��������`��<�X�ؕ�����	��u���E]��>f�@Y�m����9�މ��yA�.|�z��[�}��.����>g'�L�g�bD�xS6q��-M􉕕��2O���ńLM�+�xA�����W �;���8��<+�Y�ҟ�T���a=�e,��~�"��P���?n:v�H:L���f��N͠�Q~y��$����G��I��Ned�, ��1��Yk@0#A�i��/���ksvr���Ҍ��F�����h��be��^]�0�:�3r��B>Vj"����V��1<`���fW~�]��T�� ��I+#���㮞�j��C����#�SGRX���b,�#�	`$�� ��r�f�e���Nj���	��MJ�{�/����㶗�<��ڂ�ܷ�ʹZJ���%~(Z����H`���$$$���#�mM�ϐ��Rԏ�\�5�����]��߲�&S'&�F�q.�����|���q�!�5�ަ��2=��#c7����qT� ;�{?).���n֝Ɛ�-�ܘG�<����w��2Z<�,����ط��H-�`Cl���5��1��3���e�Ȏ7��q�����!ͅ���v�'��l>:hLٗ�Y�OL�}�G�xғG�0Ca��1fC�B0nҐ�sԟw�7T���.�&�����x�GpۦG�w����t(��a�Y����*];u�W1�K8�+s�44�ꯇn��i=;�
+�ۯ��l�Lm`���IX<�����`j�5	����ԉ\C������&��D�z�S�Me;�%�AC��:y�*z���dc�$jT�E��yJ|���y�85�tTg-cb�.��T�&?~\�����M���)�u���b�L`j�kB^^�%��I���9T����ҳ�e�o�=Y��'�����5i���a����9aERVW�oo7_`��qݨA����(�]�>;c��k#�n19U�p�0�;����KVrv��J���~�h�Z�j�9���N�g�a�}�����Bl2��N4�Ѷ�?n�u�����8���z�#s"߰.z5�e�j�:�.��l��~��ݚ��	\��J�a����̀�Wt��S��{�|����zN�c$8\� _-|j���GO�ʙ���;L�����.P+����L=mP�;�&Qg��^+����?W`[�����M(..��AU�?��|�fG�-P��.0`��o�r~��� d��e6�>x�w^䪻�bIl�Q��|�%�e���C�(	�M72ʌa�ȁr���P�$Wy.�[�k�2E�����ى�B�|To�j���˞Rw��_��+�b�����6&-�95\��d�,�	�~{�0�;F?�I	�\^�{C��Fs�i~��G���[^�\!��摵-�1|��l��C�Ŗ%���&L��u�~�$��Ur�S�Y��-{޶�sݨ�����hV2�R
�����؃>���ц�-k����6N�����{��kHeW����&�n��
��JX6C���V��D��j���uW$�����L`YZo�'Ž�d��y�w�r����4O�JBI58��WtQZ�;�/[>f��ivb���?�h[�8�Xk���R1�pv{'�VTA�nl�4�׽�J-W� ��cc�]c({�䁫E� ��������1��Qd6B�l,�ຓ���Fjj*�{�m�:�-��uU .-�B���^>�q��
��R�o'C��B��Aڡ����3]zG$4t�õ��Cd#r���qsϡ1�k��컫כ(o�re_8�E���_�c��A�*+)�F��(L�ԫ���0�o�Qv)�i �����k�Efmnn�|�t��A���fX��n-$w�:��'��P,�e�i��������v+�LI(��{�� s��w�-�A��	!����#�]T׾YU*�Ys�� Z�?}Ux$?�������[Lo\�W�L��z�ԅ�.*��?�HD�� �~gU��e����j__�6_r� �Sq���,W����8<Z	���D�b^@�����d��T�s<���K�N�%���B�Z�W���8u�hJ}�K#I��V�\N�G�B&ygl҂SM�1�"�Q;^���l�����T�Y���0�Vn��G�-ϩ(�4BJ�
�s�կ
?�[7����Rq�Yߝk���R?~V@����1�0��v+�:�u\B��Ϝ�u�ѨP��PS&!����>����^݆�������K9���u�!MV#Θ��C\o�4��@F�!�Ԛ�L_��Dy�����=��j;��ֱ�u�4)��!�,^��� �Ӣ�:��f��� K�7��~��@�� �.�.W�=i���狭ь�AY�cv�p��&~.ed٭\�z�<|)@�H &�D��yj딇F��\��dbA�l��w$�l�z�^�b���Z��iA�e6/��N�������iC��oΎ��-F)v?O'��o1�V�SI���Ԉ�&܋�#
��j��	�:�浺��f��`�b��ߘ���V.��Z �����P��L���5�d1�$٠7���*�&'����!ӄ��.���I�Sf>Q$��V���cE�?���8���B��un�U_OOO��dc��<!$_Q�;�Hz�"67���3�0�>>>0dE})�&�Fс�*z�Z,��}[��D���э�"����a0Ôt��(�\{�Bb|��~i����X,��{�K�0�>,6(~�aܢ���:����b�;������-�r�vf�PQ��[?����g��H1�	�Y������!�3�����y;2�C�.�r�K��h����&	�K8�ŀ��Kȕ��K�`F�Q��6ZH���&��-��ie-�K���e#�1^�7
.x��ƈ.�[~������f���^��Toe�3�>Y�j��At`k<,�qB���t�٥��^��r��p����櫪��>��|ɤ����;�WZ�.������:�̍���d���NO����zK�Sb�{=��1D�2��K˱��n�/�h4L�R�z�3�9�0?�B[6�]�/r�����@�̵��9��!��;ɲ3O�},�U?��&�Ɗ�����f����B���e<=�4�������z��=��3�4�����`G��T��Q��N�ݣ4������]<Z��<��@H�[ɚ%��N։5�`��w[ͤp_�ȁ�Y�N���p�B�%�)��	��/�d�[�:Ƨ�+2=�� ���%��Γ&��8D�|%Q�y��H@3��#K˨��m^�$a�j����۷�e���j� �87a�?)!f$�* u������xc�����Z*�1�Sv�_�';OsF�N,l���S�Aff&�-�>צH�"p���e���	1����cZ�8iG��X  ?���$ѥ;Gݗ�Ks���xU���h}�n���E���$�Ђ:�z�v��~�������W�H�3��>��/8���&#���qw� 8��-_�Y/Fa�7�Td\��n����l�`��ͣ��������l.��� ߘ��Y|r_���.�4�K
F=_��X'��W�3�Q� �n"�܃%!>tQ�E�l9N���F�)�/��4���M'������x�����w��x��3G�ƀ����v����y+Z ���b��k�b<�Lt��(?�5yƗˇ����/(z&s��y �ԔӨ�@�uC��F�\�����\��%Y�$I;��?5�[K<���Q��a)}����~E���}\{��=uMp���^|����-�h#u���6���q�K�Tu�{#�dJ=?a#M�4�\�&�9����O�0�܇�۹�c��Ų��R	��.ץ|�6���AP%*>OL����b�sK
��ƹJ��v��ɽ��!Gre<�vC^�����Tb��h������\|�J��H%y����j$6�Y�v���4���'j�[��` 3u��4===��F���[�+#��Ej"3�Q$U��2`$��EB�U3�ѿf[J_��m�)���eaˆ�/��fX�=�HM�0k,W�L,@6�)¿0a��Ś��9a,�z���cf�ឣ�^I�',;@-������"�A���k+
�k�`3N��IAUY
�[�\,��Q��/)V4(�ߴ�fi۞�[���
�j�Z�w��{�^��~�� ���¹��k:�`�n��9|���o�y���Ԩ�G��|��0����K��O�D�����1�P�C���H�+�T>�jE
��UM��i*�5�S�l�3\�����b����'c��!�v9�Z�A�!� ;���'������/��Ҋ�1u&]Ⱦ��Hx&�ekE��S�͞?.
ױ�	�S�� �r��~�c��C��8p��:~��P��vlk��W�����|Þ���{i���>{~f0��u�s?-��B���ϼ7���5h��@u�[`U�D��Ba2(�}�
�-�\��9SD�3CS��%�w6�t�,O�P5��s���J�{7���ŗd�}�<�� ��g��Z�Ref3�Ni���R����U�.��ʣu�8d�XzGuW w!��|��ʔ|�D4��s��!�p�N��]�;�w�k�0	�cMw�_������͈ل�O����;�����3)�qj��zH(�w�p:��ڱ���~%�r���Nmc�Rt�bL0��}�^#݃��[h�:s�'?�ԟ<��0��/>��Z�3��A)��
x ���{���y9�D.�;�X��E7߃�~��m�"Yu�q%���w�?��2]�7z��|ȏY����0�J��9���:T����s���	%���u�%&�f��I7�qO]5n�3;F'��4ߤ�w"<�k~�]kjh��}��c��G�R�p_�:E��}�����-��-\��O�x$��zc6t��#��wgR��H�Xk�F��}�0SFhEڬ�˞Ho��~�$<�L��+A�Jc�i~z�3�e�1l+��yz��Y�d"��rZ�2�1�D�z�^w�V�K����_�t� 9��1���v>�g��CC�@j��� �p3��Φ97g�:C�;�X�&��R1H	�Jk�zr���+��@����G����R������ y.eV���֟|���?��}�g/�j�m��]?���d0Fal�c��e�P#���2�vy�����v�lj�"�D8��BN$��0���l:��x�𽷊����ja�\X�|��~5��A�%��C��A�W�p��I1I��%��-�sy(J9�r ���HpB�b�K��M�[��'�ո���dwL-�ֲe�ز�];u_�*h�!�)��M~�֐tġ���+0j�U��kE��q��.��c��#�_��twu���ƸI�;��	�j*
�Θ3d�ko�Z�IZ�h!�n�H.,�Mj_o
�T�����5H��
��w{�-pq�5��o8z���_Q� �����>�x*�A�l��$��i*@ق�r�1Y�;1w0Q�j!2C!um��e���R���Y/�fd�
�Wm.�h�h���V�H��� �O��a�������TG���@X���WF\s�WL hN�G})H#��W1Z;���j|��R����)��k�JY@�7��K��pb�|;g t�9�L3�/W��g����i�Ɍk�-�9��;"Q��6��M���?3d?[0�b�0��
���`����&<O<N�ӁQ�%AĹYw���V���y6G��z'���v�hf�$Cf���l����_�����I(���g���HOҗ��3����� �����=חH�bm/i�>=yTW��p��J=��;�?8W��V��c�wq*���m��[;�Ԓ�!�)�FWA����C8���\oL�v�r��s��u*F|�=�e�8�ɮ��5�IԏQ�7#_^x��B�P�HL�#�틘fÅ6AG�<}����l� �+�����QYj3�����>�v^ߩ�ły1m8�F��Pl>;;{���	巻& ���	���X��
y~���I9�B#���bS*5��:$�p��H"���F��������ݱ���B�.͋{@}����亦�Pz#$�B��H��'ǔ�֎�?��V�.��=����]�x�(�ȴp�h��5��Y
�p1�7O�[DXxs%����9XÐ䓢ƒ�M��ߐ��3̓ѐ��Q��l�ch�}�e*�\C(
)n��a�1QL�n�d�+�`c:!��<��n�L��9��ׯ�ӻ�����	�~���&��#J�&�o/z���A"�"��ul�'cWLmJp 3],��*}D:޳�[Ik����]j����{�.��F&�=���Mf�v��vx'��)�SV���J���F�.�sM��f��0M�p2�l���p��D��]��e�:3��(ٙf���Da:7��;iQ����ِ��(��P��=K�`Z�,Q�����/���፵j���П���7�l�l�}1���ۑZ����g(��w�t����p�H��>v	

��%�£h4k�맹�N��#��#Ғ�� ��9f�X_	��`�Rwi�U�9����)mo)s51����D�&e��e��̗���U�Z\La����mq~�,n�Z�{��6�n�ǹ�[���ϙ߸�ȝ��� �n]˽����SnO���> �o�]���]���]���]���]���]���]�_�|�6������$*	=؁qA�ڽ�ՃE����S��}�(����}�鍸 �5>]O<��^9�X׷�r�Ӵ"���S�CgB�>.?\饪w��N��3T�͒OoM�%��A]/x!V����EmE������n���o�o[Ł����ԼZDD�,��� !,��c��!��%ߌЃnTgt�\l접�bB��*!ʾ�jj��?�;ܘm�����=�.FvL�O�>=7c$5����Cʣ��&������4Fy�0���q�����za�3��ɰv�Ԡ
uji�~�W�ƴ���ٞ@�y������kI٩z����T��6r��_��G��<�/�D�+�Z~����]�]�OClC�go���?}O�.��L�~6h[��ݒ4÷��Eb��ٱ�'?���E�/�ut���5����c��u?ߔGƞړ�޽{��UR���
]?U�PK`:&.Hs�~Xj��9B����@�����3�����x�Y\��]�������~��av�ҋ����&�7:z�h��߼<U΋���y���x��b�޵�\X����KW����3qu��UT򚚚���������(�bm
���n�õ��C����277��pUEⰒң��K����+�z�߃JZ-Je˖,��[R��e�E�˾d�-WFH��k��%	I�-�l1!ː��s����<���^w�|��,��}�9�s��Ae���P	q�"�Sm'�Dp׋0Aѷ�d0��V������o��AwL�C�S��?ݽ�\�2rKȤTĭE�:����A����OOO�\���b���H>��l�o߿��GO[������0�KPRR�-�ū^�RB�Zf�R���u=	�7�m"''w&if�/k�� ǈCǴ����zk>~������gҳI��A_�p�ب�Ěw��.G�����߭<+�u�����/�^�#���>�%����=������0e�9vqЏ2m�=c�NZ�5�r8@�����P�
�ء-�d0�\�GOO�R������~mӊ.���[ξ�fX[ض��J\������f-�D���� ���x�b��EN��G�^�4u�������$����<UO;�'<�70J���X{��s��vN����uҹ�
ї[H�~�ܑ詟��e�%�`�}u5��{O֩Li���*�[{K6�q��4U�W�C����*�����W��OSjB,M�[�����6*A������ס_9��)V�R�s*��ކuuu�5�5&B1Ȩ�%���Mۋ�0�4��)�K��9t��ԔQߌS	�#�f"�oF�������9���"�Z��_�1�7�S��ÿG�r3���{z�0pȦߦ�˯�x����՟��Ԥd��1ͦ\�>�[l��ۅ._IҼ~��QLLڭ[�b��s�;��<���Os�;K ���W���'?%��mZ9:�����Ν3%C��}łvN�02;Kij��!:W�4�ɹ!!!LE%�㏻	��=-�G����34�a�`7u9;�Y1�Y���-J���C�FvtD�hK�zt����e�r��a�
�9}����EuJ�9%����af�/���)��ߍ�������?_=���6^Pݘ���'�^���]����n�O\+د��s�<���+�y��G>������s�P���TEԇ��#�`\�ͮe���׻�SVj6� �Sl�̞]�|�Z #2��o_#<%"�Ã���p],��m*/��o�'�c�dÙ�
GG��ч2��^镕��϶xj�@��(����KН�8��3��TxC�NݺS�RP�{�M܄�<:Č������{�><:�d����!'���zq���L�˶~*��  ���"�ɰ "}�'Ff���|FFƜ�1Ew���ulm3.����֏������c-�̳�ۄ��^�PZ�?�x@�?�xb��]�\�KE�K�_D'��Ss(O�'U�_����2�?�IO���x=�������	U|a���#�vU��~;���o��;���f�����Ь 
Q��ݯ4�T�M�1��k��S�~�C���n�W91�)]䁮�Y�۷����`VT�O��1�r�-6 }�Q���R��,��2��1ְi+�}^U*�H��C�/^����g�G��t�;RK�%jh.�u��ۊE���*���C��o��ej�����",Gp�O=����7*�xT���xt�!�z����͹2i~�F�S&<f||�_Pp�����M^���%W�Ʌ]]�>�	��D_G,@�2�n��[���jd�E���q�/�6EP��X��:��^�3��Z2$H�UoP[�q���; "�����g�͍�2��� D��_�;���}�SQy��f8t�&��m:R��c*�f-E���u��|]Tx�KCA����!' �jk����MP������ڈ�u�o��l����|������U��Tk�+���8;
�H��\��^�s��1�YL��/��~�J�@DWb��׍���ff�k�1���]��y��mtf&77�	,#�������ʢ/!���)efh=g������u[������2��.�<���h����ľ�)���r���N@-t��w�P�X�|�����9�n�\Zm43'�v�jiY�c�(8E��� �y��`�ݡu��Vp��Z�����"�W�nQ#�cߕ�u�@��NY9Z=M�pc��vt�%X��dP�B8`����-Kkv����;<��ia���o��r��1��@Wt��s���[G|�N!߳9�ξ�<ۙ�"\'-�'T!� xu �m�v��$�hyʔ�0Q4詈��n3?5ڽ�����7n�*�gj���y��ׅ�Nx��hu���k�sKE
�.g�XB�Ɡn|s9�U�g`+���.����a�� ���ƅ	��Ww�m}���'15tW`^��}�X�}(kk7;;:ҫ�QR�K���n\;�:�F���������/�սx썅frrrܓ'�ַ�&Z�Ey�j���4W�S�������þ����/D��.�Qd ����|ɣa�-r��v��Ma�r���@̽�7Z-�7��yV毙㓼��|1�'�Sҗ�-3�=��x�����\C��߷��G_6�V`����l�9/�b�?���swͺ$
V�mK:��@(� !!�g���J"�����<�"����2Z����ILX[z���`#�`���j�>|��@4Ǽ���e��3�K+����	ɚ�>��FI����"�6/��oss�h�Wq8�xˢt���<�VN��@`�u�������f�#bbx`��>�P%�F�[�0�zu���ΐ��C��$%xfT̖�X[[㺶p���S�@\V��ֱNDWG'���>Uf*��m�\��!��[=�#.P����]��kij�x�cܹ�chȹ9cž;�S�fU�2n�~�/��˪.ʹWn�`Ƃ޼��jm��=�oz��DRaz
^&1V=��rp=2��[�<�v!�t8̼��1��n{r�}h]Ry�4����E[`��f�^��萙�L�9���^�:��][�nr���<���ﯧgf�
=�^@�u����4[��d]�Ƃ�Ү"�����M�^y�cv|r��Q8/?�?�sK~aa�2@���坌v���i�[��p�}�.��N�XM�j3c\�z\w��a�`:::�:���������tM��m�gb?�>��*��@�So��{�n5Ё/+e�+Qw�>��·���ʁ�������-���K�~���9�)N+�-{j�l���I���U����*&FF���[޲������4��@�-'�t��Y�fyKƕ�jE/(H&��֛�������f�h�8% �!����D����<o;��Fƌ�\�X�;1.N��U�,���(B��`�-���2��I��y�ec��ⱸ���#Q���!�&�(a��vaqQ4������z�G�~�omj G;�\6�D�+P"�rM�mM�v� ��޽υ�U�;���W�;��O�)�K��)|������5��X�#.� ��XD0���ã �`PX�?u�ĕ{W���rTהn4�㺶���#����^y�>�챩�F F���^��~��!N|�k���!�p+��tu�ZFF��tu55-T�D3�>6󔳅$�L�\������?����(kgi����~��~)9b�(��B�K�����\U��������\��Fط�0�����ۨq]Ŏ��D�聦-�w���<���'GA�gܥ;{z�SS���7O_�YZg���*d�ˇqW�i���*\wx�(R�>�M��4˫^'��!�����L�2oq����Ϲ�ПF�ݣ�H\GGw�����"XYi�n�u-�ބL-p�*�Ou�o�	�!,&��g{0v��j���3��!Q
�C,ӓ��X҃\��H;7D0I�&�˭b���)HcY���tP��+d�Rs�<g��w8#���R _J2J��Չx\�6��]ۖ8 m�l�j:@|���]\ǻ�S�JJw@L	�跈�A��H�8<�{�T�c���G)�-3}���Kc���͸.AQ� �wݨ���m��}v��A�rsZ�s�46^����J��|���f�++�@���Գ���PQ��~�����������E#}����AVJJ}A� 8;t�`) �E.����qܔ����?4X�d�;1q�B�٨0�b��lw��mW�|@!���o1�G-+3���h���"���,!I/^p��;�	O��51��v��zZ5�3o:�b�@,j���ڧ�&X߯�xН�*&ff{ �����Owi���K�Ʒ�mx��L�\��%�)',��������`�龜��3SSm^Ջ���,�N��:^����[��u��a�������%٩q V�J�X�>�ڗ���� ��@L�xdxi��`KT����}}}��^k<Z�ʝl`棄n�,��8:�N��Sc�?�u�	��o��n>������������6��ي9y�#��)w��r��B��~���&+Q虁�F8�_�(��wW.��RПEc�F�2j�bT�砏P�W��M���,�]�X�cg�k��r�G�=��錴B�'Z�/���Y��i�`v~���#�'��`FJ\���|vv��Jȩ�f��t~�6��G���DX:�΅�-�v~:�( �Z�ā��N�T����3%s��J�f��3�
(�2h^C�qFt#kl���-��̜N5������z���1�S��rZMU�:t�*C!�ʓ�z��ǂ�HWt5𾢒���n�2�Dg�i�R#O��>�EJ���Ci�K�m���e��։�P�ah�ro��r������u�f\����>7�SAy�����??`�� E��[�$m �i80�A�|�����;ڝ�?�����%�]cc�s�N%�}}H���Q��KӐ<�^Y�!�9UL�m�\=����QVP�dm�"���C�G�764��>���}ud:���̬,=-�羰B�C�P2�~�����D���\SRV����;�Ae!~���Z_t���:�����*��}Ŏ:��S��}�}�x���<�����{�����$i�<������8v��K��A�ij����Т������A�f���q4L�ʉ��\�_�.�32b	�����bj�]��8�4��w�V� z�����b+�sl[��@��9:�yxY{P� +�D�W�e��j��`��� B�u;:V���&����a<Y&��v�O��h~�-DA�Ģ()�����eTV�?���d�%�ŏg|'bm�.���3}%Y/��D� J�u����Z46��|(ӐH�R�ulA1(��н� ^�N�gA3mϾP�g���r~ˆ҇���5gff2��+�^�{���а9R�t�@��gt���9dl��w������'C(q��<3'g&D�Ԗ1�$���A��
dٲ�����}�ƺ�r�g�No�<9��w�m�$�Nw��K� 4���{�ߥ���J%//{223c���wSy��S�fa���'<�ݿ!����َ5�|ǁrbȭ`��oߞ��3��(q05��[��X޽gOYx7�X�)fţ�q_��\��}%���g@� l��{�I�+5�5C@L����f����o7��BPfTT`�Z�LDCd�����:��a�9!fd�����@��_�t��lȀ��&�T��ۂqK�;��#\�������;u�������-���I�%mmZ��e��N���v�����������V:�}�LU��ւ�Ru��7��Ԡ����3�a�*%` p��;&)@��?���RRlM�CVEE_{���q�4���MHA�k��y��F�����v*�V��n��k�m�m�٫i���'�JO�2Tݫ��?�=J���e���wͣ�,�E�z!c�yx6��//�j\+���]*]���DHx�XU;�Vw���W����g�\5��S����5���D��K�uE �T n�q�a�D|t7�*����R�o�e>�0��TP3H�B �{�-䒌 y������4�y%%2^�)*19X,6
���F����tHH����]Y:�z���y=��Mx� )����e��v�h�7Mtp=�M�w�V�gpJڇ�'�*5H�n���9�Y1�.$�/ !B��R�J���4�j$���{�>'��뺹�>)̦���������<��Fju"��/p8���..�����H��[���7�AYlq�6JW�	��������>�V�j���z���V�
�I��v������q��||m�3}@E�M9�����L���bd��A���Y`���e?�Yii=jjjBO��:�2}{�<��n�������[��-�	�BLM��@�`��Y�2`�qq��Ӏ{ cs�?�`�����5��h�2�l�[�.{�O9���AAA\ǖM�km���3[6ɑ ��-,,��-,,0������c�~=B�.~�\l�r7��+�ˁ�PJ�R�`�6=ݎ��q��4�ǆ�(���Ye��}��Gd%+�w�v�!���?�}U!=ݏ�!J�-�wn��+)��WS%d��^
�ۑ|��=oԭ�t:�Z\𲷲zWby�.�8یG���m����������t@���,���(�g�Tf(O�<���rGo�� �Xp���)�����/�A�֕�����Wa"�}K�����#.=�E�%���?f-��R�u���>d�_jS.�,��{VnU_Ymhn��j8ߣ��(�l Ef?^�m�KK��/]����˶������ܹ����%K��	ʱɫ�繒��� � �!��h�U4���a),tc���2�R�������u� fɱmx1��� �+��@c(��ڟ�]�G<�K�A�l����V���(Kxߑ;�hJ��T(�ر/���}{���#�hJ���!��!�W���,�3�����J���oƺm\o��#!�ϻ%��V*��FB9��(f�Z���֕g^�\1�D�� �|�v3��C�=	,c�tX-ԁ��SP�j�
<�s�G7�:::7.��3�lw�a
?��u���t�I~�ϋ�@ׯ�	�p)Cw�\�bŷ
�:���i4\����S�L�����7�m�I~)���P��$AQپ��mhh����Hc�����wL?Ozݸ�
�#�A�2T��de=����]��[����T<�ܴ�]��[�>d�AK��'��z"-#uW���"e
?{��? ����x�"�͡U(A�T����������6�C[XE8�X�R2�TQ����ܺM,6�Ύi9�h�10�s��.�n���׮�|i���+#Sfz����EH㕡@�T�TR\�{2���_ܴ���]����{�ǧ��x�������SSZ�	���A�����Ɵ�b�S��߽zS^E����{���v�O�$>�&e�HC��F�� ��a�~C�gh&I� ���8X��_y�S�)*h-#�Ɛ�,���B�)~�B����_��H�BҞ�6����E
��
���A�gfj���oqc�S3 b�6��(�25��H� D+�@�Mjk����_�Ʒ�c"PQ�<g���44���732*{>�/�(d^�}��rJ:�>J=����ֶ]�0؇OX�����P�y�����Z���t߀�\TH�cnn�DK<�!'��r���7�S�1L��q���ݒ�-�Z;Tm�����=�o�7��E"䙱13��0����J�� ��������IOI�^<Q\M�K*~�;{������oz�����K� �_=O��m�(&�ދ���D1.� ���7��hq����4��!��Qd"�l���o���`�Rs)3�-v�G���}�_H;c����������j��\f^^k{9~d����^>^=�cu��9�B���vԘ;p7�ʲ`�X �܏Z���-��<��;���߇��9�20`�q��^��=�G�[Z[K�����sXԋ��h����P{9��d�xbX�(rDjj��)M�J�B+��IvW/�\�����Ȟ���>`�M����_	�НW3�j�YRҽ��Ъ��Uo��,., ��_e���v�
��k{�ɹZ����
C(v��a����k&^����_�ӿ�ʝ�y�f��<�r�p3�p��9NDs�(m�L��x�R��Q5k�v��c��
�;��*d�2Й��]\~ĵ�k�
���QX���߫���3X�O}���UC6m6JW�9U-ĂO���랬���۷o≈Q��L��������>�����?�>����,_���̬�y�w�%��Fm�;��s�~M���,�������{�8ǥ>��pif�f%�)��Z�������@[��L�v��a�55C1�e,��M�5;�H�\���!����=[��<��HƂ2w�u����� S����Vﰐڹ�z�۷�	��oa�8��S�U\)�n��=��� � ƫ��=�Ɩ���%(~����e�����ZW4}������{Z��g��[�ܚҟ�݂�j�iz��J�=ܿ_����湴�4@��9M����Z`��8�=�
� �m+ﯻ��4���(�DN�NBZ$X�v�:e��P9}�5-M����?����nnVZC��j?	�������rPx�kB#Obae.�?�ZGf)7�~����j��zwJ�i���F���V�Y ��̯v7�� .}�"����Y�N.ڢj��YR驧�!��F���x�<�<�⒒Y��]���g�[�����Ӕ�4��	�����t͵����	���]��UX�f4CV-�\��UT\l��-�[r���{YTbm��;�H��{�Bo}}=�y�W�$������Rn�V���@���R	����v�fr�������y��싅|D@�����/B��� `]	�u���
��C��.
�f��WY�P�޿��L�=�A��,�G�y���&(�����"9��b�/\�g�Π=w���'��T�o���l�q8$	M:>^��>W�Q��(��'j�Ѳ���s�t��5UM��y��@�W�,R.��!�?wtt�%�;9!�/H���/��F�����Z��Z���YY��>>>����V*[UC��-�A
�O��4���VbA�����������<����B�=�=�����E�h����ۜ�֦EOOo4�f�!�/�k^�)Q�sl�N�P��)���$�D
ư���*�C#`�`�B��B/~Hַj0ky���ʉc��pG�I'<[��u��R�[G+E�4�[J����M4CR$���,wbb"K���Ȉe�ͩ��U�к$P��;'àҗO>�C��.��fn�
M�����������:��@�`!��t����5Z��$�N�%���׻��D
��͖)�'�.�r�+C�Y�,ʟ��j�v}�[5�?����O{|�����pׇ��A��"��t��_a4��՘��3b�b��3RR�ɀ ���p�v�w��%9H�̝A�M�W�U��ds���G��l�΂�F�%���_/^'*ބ����Ń�v����1+Q�S�9L^�����')���N��w}n~��8I\L��ǡQA\H��
Ph�����^�B򉪹� #���8�,��z�bT<��A�o�en���7���LVq���UB�p��0�,�30�k����A3��鞨��� {�ݥ}��j���-䏐v�t�U��B�a`.���
�TT�1wi���r�%555��r�x \�.9t���� j�m4Ui@��6lQ][�Y�!�s�FV^u&��ҧ͆��E�S<C҅d�f{�,עq�Od�S�gTl�W�?��j����K�0���
�L�t��-�P0�8���stLX	����g������"d�����:��T�5�u� ����a��i֢��o����������NR�1�/��da��~5��˙:ۜ�O�ӈ�_��n݂J��K�î'2G���E���K��"��h8�V�	5�H$���d��}�"V�*."b���? �"53����������G�S؅<�I�=X�in��/,�Z1P�0m�Vڰ[�O����9|������Q��r������`�I�܊���� :*?�K���f��sC�k�+�QW�ڒ�]�����>�гM�7����:����Yۏny�0Y�V\,�%ťfpR�)����� ��O�@�ܦ��3��������
R$��������b�O+T��Ҷ�cA�Ν�]jSv���dC�RTG�Z�$���̂�O~`<���i�b"�H	��Y�����������!� � �ߋ��Qd}����0��i``��+@ϠL׉8LQ@'|��Y,��ݽ��j��u�LZ���% ����ɪ!<�*�Ӎ�%����Gp8�_[��_�.��R�G0	�G�à��H�t�}���&5������S-��оڦ���ؗ���grhӶ#�j��>�����#.h^=��������]��#�����m�"��3��kg�>�����0\���HS������OVy��SaIԆ���9���YT���{���͉qځb<%Ƭ=C'�!����#5�	�����?Y4��Lbecs$Ty͙���7w����'��>��_�<����t�^yE��)�a��������'?�2�]���B�Ho�<؂�,�B��x��,�\�]�����)�J�F�*�6U��1ƕ;����WT��c����r�R��n��Ο� (Q�w�PЦH))��*䋎������s�r+O�/. _�:_�j�v����K�|�W�1��>b�
�qb�$Fw.^± gel�e����/[�\��F���z.&��顗K��;��XE�_����붶��ǡ�j����O�4M-���g�+s�g��#1+3�t�Y�t�/M�T��e��n�����@�:V��ˤ��oYbՏ�IGY�
G����6�'�����(E8(>��z/
&�, �:.>ޚ%D�Jߑ.ߴ�#u
�I/�!v��=�$�/�����"��Q��,�TU?��vX]]-&|���0��,<@�#��H�Ñ����_�'G���27Ot��2<���u�O~���"KrJZ'G_�m>[\Jʖ,y���ޖ�����䱃��1��ƴ��9����?.���c�U3��i��bT�̜��E3x�vF8��arವ܉%R~ܥ��|s���6�!G��߅6�
@�j�\*vo^w�v)�&	_�:$vP��ħ��N���Ҟ�Avvvߩ���?��-�	Pۀ2:� ԉ\3M|�$��NC I���/��sE(���0�_���k�!yD�I!���=�f�����=T�#����o��+*��Dk[h�����ݧ4��ۡ�f[��bç��P�-v������F�	v��k-�eN}�<v����!z����w}u�qF�cSS�QwS���D�smm��V��k#�����-��w#A[�������0N��2PT�T�/���7���k3@���&$��1AY�ĴŦf$�������C<N~�듙���iV�x�����;U�f�T�D$�U�/_���s�[Ip�Փ�*��zu���.by�4B�^2�}����9��<��@9��ě�r䦧�ǈ�6�I���T�OyN�8�KH����8���`��3j:�
��S��r #�F>=xo�]��"jn����ts{MW���%����Gmx =��f(��o������9D���4m>��{!�k��>y�)ƚ�Q��q�W��X�����?���ӝ���g^9HKy}�j�?���\�avW���\�cb�z�h�9�\(�2���ə;���T� �����E@�^�~?��+__I�p$�h�F��y�g��,G8�]p��!�L��k�E��ꑮ7}�97(��j���ŗX�e�c������dVR�e���ҝ:K����yo����׹}r�������%���E1��X�ll��~~4~&8�XzMM`������٩�@)op��
tIJC� �m�l%ZYIu��۷���1v��}���O,=0_{۵eO<.�.t/�+��+ ���A�&�u��D��w���A\�M �Q���7WeC�����Aν/��a@9p�u�^zz�����Mn�ޯz�\'���n�{��.?�i���U���ZP%�rFL�^,�T_W�ef&����X�����L�����}	�}d1		��z�8H��AԶ�K��8K�	i�*�g�p�6_��x?��*lT�s��9��..5$$�af�����K@Zʫ5��,������`
�S+F=�qXY�k��u��������o�m)R)�����7{��U�S�qK�]�;M�6/�j5���ps
op����
{���I������ߜ?y�����ey芠���
��mZ{���x70ٳ���y��l�n���k,!���s�va ���?ѫ8��fh0N+���I (�{�p�=�D��`��H` (̽ T ���zތ�S��쩙_K�=`W�f�}��c7��8������?�����>�4�/^�lb�`ge-�3�{��'%@)��T.�f dy--�$޼�ǉ�bvV�Fc>ie��w2����h~�p�>?�пk]s2`�̬��U+#u��Z-����Zv2�Q�	S[�|8�j�0Gt��WyWGG!o챩e�U�lu��.������'�Ur�-v�#['�ޤ$%�Y�N�]��c���۬3�h�.&�W��_m�j����(u�/�7#S�`(�н��U{�:�Q����i�P&���c�M�ITMh��ɢ�,Zd�ZIQ�Y����ՏN;C��Ҙ�ܨ��k����f��KK��װ���=�9in��0��}O��9���.��BOf	9m����g�L�X��Q��~W���X
X�b��)��RCP
��T/k�^y��P�=����}Pk�6�R,iؑ���>���,p}Ui���, ��G�-�0��Ra�˗/C�q�������iX�RWq�G�}&��T�V��aj�sWɋ����~����;���5��T�$��##�U�ي�Y�'!��d�}Tk��7���g��mȤ���ڮ_`������]�����)������#w5{��3��}o�/~����{��{,`w[d�R�����q�ǒ���H��6�w��%/��犖[N�3����>@���O9�gC؜x�g(x���&�MO�n��PJ؝q�{<xp���$ǡ�A�%�*v�~�Y���ʟ�%�_�0-���36��u�m�7����P�������Hh��h<�_^%��=�6�?=�:8���k�s�hXJJ�7�Q#�׿̲��^���z�Md��Kn�&�������U�������g>��̣����9��e�LLL
���z͚���t���<2�䵸���n�7B�����S�7W:����[/�p�8��Bǆ��oWcH���|��U��}3������νa�9����1��C���Չ&���ש%4�����V�Z���%�����4�M|���\Rc�d��>55�Қ����ݭbĖ�;c�Ɂ|s~�U����Z"�٤�X�o)��ײ�gj(}5��9_�|9��mb��WxfJ6�nk{�6ݎ�-�����;�R��7�afy���o] �Β�~�{4�O>Q�#3�#xz�]�ЋU��n2k�2^'ńu�nߒ��Yo\NQu�[:[Nx1�>�챾��8���)��m{t�� �����L����-)�t���<"�{q�BD��a�s`�N��e�z�w�S>{*b�0�IQ�y��3����슌eԙ��|ك$��y�{Jȭ�-,��s~w]��Q���,6n�؛��Y�jU3�[�M~�.ذ�tBK+�^���iwq��oqxUD�q����^.jwz��u����D}�}3(HM��x?%Ȕ����$�0Qf�T�6�{N�:5oH4H�)��{�.<8Lt`g*�i�,1�3�z�J��Wџ������G������.��=��OL2�<M+�ߘWP����d�?��!gZ�w_�~��t��T�-+d�����]9{�) ]�R\�0�.=?�X��E�j��Yma�ۑ��	����j|"�����F�_e���Lkb�8���1� �x�R����ڸ���-�T6���+�^�u����!�ܹ�޵�����v!%��#�K�o��/�o�&�� GRA�~ҿ��[;�[�����
�
�L0���d~��Uua����`S{{�6�2�-����6��l	��;`�f`J9d��}C�;J��&�F�`b�@���K"�5�v�p��%y��]��-�XU__�e�v����1��ͫ�-o�;��6�.f�� 0a�#O�t��u�U��X[���h�.�#OD5x���#i���Tt=l�+^���5k��G��R�a����h���<첷ظ�,�C,��>�A���0�����v�v�S����Rm������UKˤ�"N��knRo�*���l�K�y�(����s��f�x���4�z.A�
��`�2�G��Eq��o�vuu]6�Lw*a#�%��k�w���E������gu<f�Aa��-AMCÙS��\;^�Sp�z�8W5h���36�M����5\� �%��6gT�D[���Feaᘻ��^�`��yӏo�Ὓ�v>���{��8g�7SO����@�V,���%�W~x�^FFF{������cfڔ9�@p��������UEE±g�D�.������Ӻk��[�f@\;{���p9��8潘m������+��H���A$`���lvt��/�ޏ޸9)3������q��Ys�zZ1�t8��#���3�~}��DeIߒSr7y�Iug�����eS7�7��w���B��D�k�������"5p�ܚ{!��W�Wj8mZ�	z�I:���'��5Rr)Us�ί-6�il
�w�t�e[ll�ݻ����o,4�I�r�3�G�|Ōs�31U1��� ����9]ōM�3#3��/x��.'˳�]�>��]�)�iF9�n���[�x|`W8f�rI_����{��9-#��&�h.q�/[���B+������)�R�����Cr��OE��k�'�]_�����״���4��>Vn�Ft�m��V�E�7~������6sw�&���H:��{� ��}��ț���H*���˗��k�(�6j@��n���y���Q����*���uE�%�z��3�f�?����־���3T��ᗽ$^b�) _s莗�D�l��y�t-��B#�
�ے���ծ���t���y� �ے���'ܷy擺ES,�����rF��Kۅ�!�m���9gzI��Clll�_Q<�Wg�j���ӛ�.�<0P=���u�]��r���a���Sp��1]���Z�Кڔ���Z��۴�߶����Zt�)G?����W�����"�Y�������z�
cQ3��%�)j$�}�בz�5��5� �H��(�N(�����������Bss3x֩$��V*i���U��<CԦ����������xR��i�˱g����홗ް{� ��$Mg��ɔ���υpǜ�z�z������Z�`��|���L���!š��!���u(޹L�4F���c�.ԗ�ڈ}�ė ���W�d�����([�_�zs�_�)8l.p���WQZʲ����nhb�~����������{6����� ��n������h�c?SP#m3��\�K>��� S���S�[Z�;:t�y���t4����D ^�oi
ۧ���<�f<���i�[g�6c�J՜��&9:���S�_ꢍK�&�[���ϊ�>�Ȯ�_S��4�Rc5 4�Ibb�^H������}3�2P'T������	~�A�j�Ο\�s�h!D�R=#e�S<�?�7�OU�aF�R�54��2&�7l�׼ߡӟxs��a3��#� ��^XH��!�2����qo_ѥ�Q�sJ#0����������C��?��S�5�j�G�$�?��y���H;�0�@U5�Ø�Q�D1"��V��	i��P	��5���Bϡ���B�5k�7�;2N�����֋�S�@��R��{�>�8_�����Σ?��>D/����79�^�&��x��Q��ov����ѱ��K]f0����;z���ޑH���<�J@��~
#c�VM�.$����jl����6�rU���NÃ:U�Y�n�%�[>}��U�b�T�N������,��!�5���%�������]���v�'���<�^UXK���j5��� �ba}v�:%n�@�z|��'Q�X"Ba�����`jj�k׸��
��@Cw�Z�D��,�/�7d����(���/�����V>�������T�޷"�� g�^����9������3��7!�����9
��6����5���gm�@�=�_��_�L%R��4v�#ú��F�v� �ɚ�Hm�s6�A�-�q��|������1G#Χ�/�����fo@���Qs�
�V�E��`N�C�4.Ҵ�Rr������l�R�Yl./,�5x�}l��Q�	�&䣚δ�F��X���T���É��A��U+ğ��?C�6�0Q�Y"S��W'#sc�c�"����w�ȸQ�%ǻ�c*��ǈ������"������Γ�7���#���"�~�x>�[gv��o�ҍ{f!��7d���!/$k��Kg �k�4⨮炔�z�Ib�"He�?�;5�(
�\�b@{\|۾�0����VN��mtp�p�+�0f�X�F�B$Kxå�#�R���54 7.�����(i����R�a��v7q���N�7�3�	'��ܿ�3���mvd:����F���bu��km)�ڜ�/�"I����:�JUA��<"�n����EE����Kg>~��Ms�H��m_�IS�R�N�����[Zb�Z���kn%���)b�f���-���w����^���h��J�³j[
�e�vG$ԏKgd7�/u�� i��/6:�w=+r�Ntέ$����-��VƈF�P �����#�s�攳:/Ǎt�q�F�Zy4� m�{����{�X�B����U�G9!�R�8��A����Lx�FoT.������J����B`v�~SF�$�2�0�
�����>�N�iص'淹�;�?�=<�$��/%�8�^�5���p�l�!��N��"i�)"��[(�R�F����1<0�p�I�#�!F�D�s��j[q�U��l@��U�S���e}���zT=��x��R�W&
i��l��d�c!��l��H��ٽ7�
�����n|�QPa���m^A�M��~s,�K�>d�E��G.�QُC�&����h��Q�.{ǎ�����z�x~�#xx�EGY����� �iϊ�����\\@#"�͖�>8ȸ�������<�����}1�j�5��C��،��`�X��v��Qڲ�J`X!�����{����T*R�m�I*7�iT����鷟>����'7���ݒٷ��Ș�e֣1l�&�6[�;u#�!�s��n��)�灆EGG�����~���Kx�o��6N��ߒ��mBڿ�g�M��T�_:>>��3V�Y�i�*4kԱ_b\�r
����m?T����;��L�@j��!26]�2�E���O�Q�B�8b<��vl�J�|A�u�՗{�X�u���:�rG�{ն��*��c�&�H���ze\uh�q����/������06b�1}����<�3��8S�p[�mx00���D� 0���E��;���\��bbt�7�KSs�Xl�ۥ��?\���� MM��-����&9���.�m�
�i��/���҃+����Prl������NE�ݳ�]~W�i���`�fGN���]*�%�Ner1���J�xK�X/�{���t��q�g���g�6�VoYuvK6I�߿q!��ͦrR��?�����'rKF��!�2F����5N��s���<Z�N^��/�<2�G�.X���P���˙��Vǵ�K��Ϗ�Ќ븄�`Ѡ,i%���f΁� ��,6��R��W&�Ŕ�E�����&'�-*^��*U.�/���G�H��:z:c�����v�F��r��R�M�v�N�����w����Db�� :��su R�ơ�'�K��E��Iu����,�~�P&��-�X�o�<�&h��&�;]+���u�H��<��e|�8Ƴ���$N* �s���j9�~����M��y�{ґ�_�����_.Y�O��O��1�ׁ�M����?�m�y��t<�)tڍ l?�X6�P6۽i��e�#�o�)3!�W��a��V�M�D��)Rq��ڟj\6-�?�V��L}��dϤo(rt.3�������:���ЯM;��p�������9����`Wd��at�X����;&4�-�Lj*;�h�}�;����O�_�6�h|�b��W���`�����Դ4eoS�!jb�"�ɟfs>Up����[�SV��@n���2�8���(�^�o�3g�@a��t��u4D^�Y?�O	Ϗ� ��RzD�~n�f)��W&��ƪ����Ǻ{�Z�DCQY�����GE$#��]���<���d����P��d'�{�����>���}^�筗�=��u��{�s�<س&s�z@�q�`AO�/�:����#����ƾ1l��une璻c��+jv��ݹv��{�ǖ:�I�Tc�"���{��.�k�*G*G*6Fn̸���(f��G����4�1@��I?�kT����uZ	|-0'��9�m|�a��ᢦ�|�#r�#�"C-�D��3�0Y4��`��J����\�g�z<\uw���%����M���W��ܙެ&�p����9�ğ1^+/2��b�]�����&�br���m t>�C /n��a��t����釂��W�sH1��mee�����k������"k�b��&��BL)I�'��k��b��Yhц�o'�b"����\������qhB�J��a@�XBn�j�T�J񄔮u�����/$�޺���(����"�pL�/�Vi�$"obգL&������70�c9o?E�t<��D��{y�-�_2B�+A��4*	�M5!U��U�����jf���/Rc�A1Ld�"X"|��#���~5�c��u"=!�O(����]���}��\T�
��N$q^&��E�%�
#���\̨2��C�1u�NJ�{�n�d�.��^�@����}%�g�^��~&� !�;V�bG�0LѻW�C�KHSj������~ʯ,orA)��0��þ�$���	�B;��N�G�~'��d�aL{�Hq�ڹ,���P�+�j�j.��R���?�;.&���RІ���۷yLg��U(5�*n������3��':��
a�ݸt�3�Ԟd�&�#�b�E>���e����v�B!`�%(�r/���r�3;�nr���c��$!�:p?ӗF~�=>>���U�)�`��I��~������w-����}9pᗡ��:��EMo���'3*N�=A����� ��"�s��&��r��h�'$�Ø1�V�	�ʄJP��ޚ���'(�+o�1P���pc㕦*?�m���X}[����| v�O��&�Ҿ^���^�Y�t\nb-xlw�p�����􍳩=�ō�V������	J��Q����U�<H���,*�`�2���}�>�&<�:/8�Q`��s܂�z%o�N��R�b��ЫD���7�a<���g���#���bf�����|:�����YEL.��(��~��,��fΓ=�.�b���Ƌ�����)	n��M�(�HŠ�ld?5�bl}cl�!שR$���}�Н�^��Nn�[+!��LxZ}_�~�U��U�]'Q�ƣ'�]QϢuP||S����p�)�)(y��(x_�- 3�n9�y;b�s��0������G��*䑆�4��\��y��\�_�xlv߉p̣�bc���ӧ+���y̤#��(���3	�oҫV7�׸�[ösnQ�b���֭�YY�LŠ�1�KX�8~���,����Ezkn���_Z��O�/��3�(���z\C;��ܱ0�sI�#E�	��V�wh�B9��?&��tP0�?�	yL��ɉ&6�Z3�lrV�����W��e$�>�*�sg?������پ脱�#G6��u��e${IV�֐�3��i|��Ȫ�n���;%Lv�h\�=2���{�i~�$����=��T�[q=�J9JW��:,r)�˹���:�&EF	vs���Osw�\�mK~�d�On0T)�<�%���0<6O���c�� f*I���mL{+&������S�LcI?������	jq�nQ�%��#�l���]�d����ܘ�UX�u�}�����;
�O�n�QN[����?7U1�T��D0ڨUp0�Q�P`�S�ۛo2�{,МH;����ų���I�6�Ԅ�X���]k�����I�	$x�|%}�ki�d� &{/Su'P�ѯ�+_-˶�B�����r)ʁ�$9w*��c򟝜h���J��)��-����ZL.7�j��5.6���zJƝ��|��9)��	�D�O�XV��vb����'�YZ�Qn�A3��GOL���^J	?�m��y���ى%�k����B����Ŷ�'�ʛL[�nَ%�Yc\���k�$�N�C��En�oR��'���6���4��F��xWP
���x*�RMY�5Q�w))!ۦ�|��V���*�cOp$�[{go�N@�M{�O�؎�ib��W�Dj9�wG�1b=/qs�;�u(���\�~����GOH�8�t�?��QI�- k}��D��Tl�$�kMM)��W���7�`ҟak�ZR��[	��qf�����4`������X�6����t��~������H����f����j%н�=ֽ�l���}�8Ĳ���O��!���m-���*�����(Xz}L���!��ర�RK0���l�R��_ܪ�Qq�LPW�}n6r*o�+���g`����>�m�`�iI;V��|�>��.��S��66�O����+�^���]��e������p�-�m�	������lł���0���(����$� TE<ҜM�S��c��n��x���%.$��ؕ}l�È#��mD�ƆômO❰
���hZ���jٳ�9&}WD��B����{m�����HF�?l_�_p�'��ݓ��x�����{|d�֋��Qу��n������t?V�Qa� __�@;K�q��[�K8���΢��ע�)���A�j�� ڮ���z;!8*�9�͔��	�t�z��S[>l�ā��tO&��:�j�F�OW����N��Z�u�E�싷
{�Q��� V5���m7Wc��<�n�Q�o$�����������ژ�нIu1*.ȋ0 ���b�S�����B����Ln��<̟�s�C¸�lCG�I�ku�洴����b �p�&����]� �R��H�:o��:�mM��?G���P�:C[6`������\�V0�)��BC]]����W0�`2��p%��b6�L%��
U7尛k�G��X#�݇n5�WP�]�^��Oe��hW1�TQ������ŋ�*���ϻ6p����Og�h�]�jZО�(��{��^��nQ{$�<}�RKӜ��8��-~�Hs%@�" �؀ln~��_�i�NUUn��O#蔖�q�E���\Ksc����������R;��1�\��zaL��yN�\��T:�}�^F���Ke0L��qs}8�xgC�R���x+�Q�>�޼M>X��^���ܖ��Ϲ��bA%�mP�	���R�����kZ��>��r�EtB�%�cS��łI�k隉��}u������s������4.J��!5zj�mjҚ8FXoʯ�?_8{���BI�rd�}�e�눛��֒���5�,� ��~7ġ�p���'B#E�ï�H
%�N)7{sd�t�!~҄�mNcT�d�ׇ���r�⪪�ህ��0���N�������'�m��S���檻0Ҡ� �1�_e��@	���6�~@]�'���`�/�����[v�~OJN6��n���m��������U��Q����K�t�ä��g՞��,��>ϡ�[�ՙ�+�)��u��Zƛ�!�>���

����0�#rl�O'�%6=��k-��ln1D��wߏ�����^�Ȥ�n6GV�0.D���k�g��d�f%�kn6����|�A����;x~��BT����+��f���Y��z�x��k�G�̎�w�n+��ɰ��-Mr�ΐ^�u��VcDA�����/Z�2�A�Ң�_�SGL{엚rz�f�����5ʽ��lOz�^�R������묯����w��yf���;�.�} I>���۳����-,,��Dh�/4�o�#t�7|t�H<�j��O	[��fZ�..��btX�j�d��9G�i�����ӿ=�j�[���)�������W���6�ʷ7H<3RSSWF g[[[%^�w�B(u�H�et3a
����ʛo�x-�`�ky�i��E,��xE�UsyqR��X����.��t��ǭ�x-�nt�fK *6�j� ��CFgg�>q�����_��*���'1��{<���κS��8.��RZx)H� m
��Uf��^��H\�z�|�n^RW5���Cp��A�����,�1^rn�����o=�v\���<��Oe����dCL��U�|��N���c��D�BA�����Y�[��A�V�Bڷ����������_�Hf�ɜ��M�b�BHn��oq������9��`Ŝ���QF��y2��3=�~�3��z�,��$�s��w���I]�l��22<,_�X�˥ߨ�Ǩp�z2���VKCg�����.¡|��s���c��y�I,�8:F����u�(iX���2�2=���CH3�M� k
߈��kj��EU9R`��='y�����P��e���Q������S��C"�÷pm��"��)��^�E��XÈL����xY{&�z(��/�@�r�ѢH���C׽GQ燙���yi瀋�֬Aq��9��e���<�}@�i}�>�[�ī��� ������de�MjK3�N ���P�7��P���`��U��x���N�_�UD��jj����������Ϝ/��	7j�G^���.�2,b�2�d�kPlJolL���mL�����ws>v
b0gz~I#K@�ҋ-j���nQ/<=�[f]��t��)e#tF��r�|9�1i7_�Y\�=0�aDm�p�Ս��M�NT�k�E+��-�x���t�{�/}���������B��':�,i�LqQ��G�H���h�2��� �;H�8L�J��
8���{Lb�������}�\ٝݍ-'~r���z��◚�X/��1o���F�ψ{}^�磍�����!�I����cű
&��?=A-�7��X��x!����)���Y�ېfA���D푙?i�;����;!��Jm�
9�jҊv{�lA��bjtp߂�xC9��kW�lG���K}�d�H��Ԃ� �9��ѣ���	�܇e�,�t����F'K-��22�ҟ]W����>��0ʕ�)�M���B_>�B���lÈ��������%���e�a����N�.��:���𝞼�W�|�[��xRfY�e��_�b �s�z���|�D�gk�	���Ap��]���Bu�����|חEC`K�Ս͌Z�����;�jq�hq�z$�*�4fZ�G�2�2ii�Ŋ����#/�\&͝58/^<���|y/_�W���m8�eG8u������,��kY�2:�(My���4��v�$͸{�������-`�T�u�/�\юl� �}@�az	��������xr.+�ȡo[2U����}R���A��!D&�!z^�Oܛʓ�ʊ���q�̐Ʃ���'����7�wVc�5�y\�m|��V�Q�i e��/Pj��x������t���C7ϡ%�O�;����Q��!�kb��a��+���mo�F�7\~JF� �U�=I�_���/�&���A�����`��?\6޼O�o���u�ten�Ҏ �+����]��`���.Z|�/b]{���э�]�K�~��i�_��o��51��*��>�6�O��q&��L��>T �a����HP�sB�������]v�s�ϟÚS�'-�;�'U�:F�I*�����~������z�B\����J�ka[����!�[��D-�Ȅ }�l����{r\�7[u���Ð�!�q)Nx�|*'9Q�8n#���%$�_k�#�5�~�"(FE�\n:�(}s�s�!3t�1^뽘�)J�ii��Z��9Q��*FX(:��,��x��2�	22�򊯺\f��_Q��0Y�P�2|���-<��R6�S 2b��֊�|U��V�2��2��%�*p�Ĳ�afǢ��� ���CCC���5��Q~�)%�u��tL^��<���x�`6 %�k+�-�,-͕�jLx�x<%O{�w?��G�$��7�����T�R�ٛ�t�Q5�,S�uKV��i��bJ��Q�6E ����� ��m���B'Pn��)��3H���@@�>|��׶Y�.���^����گ�{MkX�=�{�w,ɛ��	�ex|�zy6�DA3٧m4�R0��F���FohJ�Jjƶ���ӟ!��������ߗ|����0��->+hH����)��8�k�KY+��0J�d��3>���O�t%��j?C�"�7m?}�򌁟_�\�րә7�Vj��������T�k��>x~7���Nx��0R��.���Ӊ��ۅJ��/} wtToK<`?�a���Ą״�m:����yMW�Ź� ���������9#~����ڴ7R��c)�����\�垐5�Q���Y��LNJ��ح$;�/�>Ik�� c	���F2��������C��l�lٹ��~-�G�Vx�Ix{M�^��s\�_��r�U���66|�Ϋ������}�:����dLC�igZn	)�N�2�s�������)��4��e0�d���6;�k�_����0����!��k�F���1��k���H�����R�N��f�


�����K�[K����
�s��˟�
`��<��m
�a^�j�PҠ3��~�t��ŋ�*��� h�Z�����Ͳ�z�AB�CP�� �=�т%+S����-3xN���l~�X6\ ���x�Y���6�I0�La�7��Db�;�k�W�zVYlw*����33�رU��H0t)-��s��|���2�Tx����詐� ���7�r��Ӿ��Y�1���~�eo˰���!���|�d-�څ4Y蝑��/�JÉ��\VV��xS�m���4�D�~�Dm��>��n�#3_8k�C�."X ��A��erq�ˬ�e�׉$�KN���۸o�1UY:[���5��~M��;O�������M�ƻ���=j7�

��{0�o�~!�-,I��"G*ʇ�/_��:�`"�kA��CJ�!d��?�15�i��@yTw~NJJ╫:-C7���~Bk&�Ğ����4�g�(�d�OOg��ED��V���4�Ʌ�)_�`� Θ�dm�m���GǙW���T�����2�MH�H������9����7G�7p�%���B������ƛH�0�eZ����*>���[nl>'�`�=0��39"����StE�Ϭۢ�SC��&�V�;��+:K��^��sb���mug���,-HK�k_T6�jA^n.{o�R~ ���khی}n�B�˴���,�"}�>�f ������>/��N0���R�cM�����c��n���qcY�яQ�G������4����]|�>i5�^�;Ӏ�z��q8���&�:�i<1� �㼸�?ߵIƋ�Ĕ�g	�)^8n�l���^-�Y��Y��#O7�I3��{أ��ivc}�x�b�<�5H���e�2d��+3�>�2�i<�@]��Xx*�_��ml�	9��m�-�$9�� _�׽5�����i��[L�MM�7�
�,��'�8��򉗻�J`qkE(4����d�Ӄ���v�w��S�=�6c�/��5�m��b��2;<�Fj�J|0]v��V�~�w���Z4�6d�T:�E.^ϼ��]F-����3ގB�u�q��V���#��駪q�HI+~�~�R���а�k�~p�~����qO�!ćЇ/�=��&.��̓9Ξu���#Z XS�аF����Z2z�9T��[[_�T�۽ F�2����3�OyR���ػ�zYd[o�9@����%o���r��z��oj�:?
�O��3���A�k����y��K��^c��q�3ޔfff���u&�����ze���/��8����F�0�wIIb)-k[m�s��S��s�]��\x=��?y�!�̵���D��2����?{M~��΁Q��2�<�ldhh���|�P:�aK�kF�Ǔ"4>���)�;��Jp��kM\��B�U8n�:|)эibjs��dz8��jG�qAw�M-Z���a|t��6�s���i��|�������2{b�Y>ټ�n����fJs�l<es,%�~�)���q���=܆_ѝW�)��;���x�������
��{�����ɺ�󩏭Oݣ��+;�՞�ͥ�ر[��;D�ƫ��o3G(�	�T�AAA&FƬь��KBڻJ�PÑĴ��QF둲��tQ���K%���T#q5w�Y�f��L���`֜���$հ��&�����k)�S�˵w�5��)���D����Z��U'���4��y�����19%���$�<☼�˚yzo&�yϐ���o���P�~�}��r|�����"�6P�]�*#{%�ޢ�Y��)=���#.�������=+^�l�2��Y����U�9J�Ϙu�A(�h`��:�1� Ռ�u��X>|�6�cF��_}�%w�����,h�� �g��oSS9������%��!ܑ!�r��KI^M7��������)�i�H�5��Y7:nv<~(ZL���¾}����[Zp7��D_�=nue�9���ɀ4>��c:p>W#k�Zm�,(5��3��.ԙ}fE���P�[���ʁu�^:ʒtGv
#R2�����6<6w�l��@��;l���Dl�L�eF��G3U�HO�8��Z	�Y�}���ų�	��8=���K[ߠ�k2�&�s�jVϵ���m���E��˗�����u�R��N��C]'�,��CQU��%S	��a;�� �W`:^��L:ka��+��s�!!-�h~��Ӛ�'|�L�5��l48l�?�Q�U��j��yuę�&�>�Ȣ:lN�YV!R����7~u������n#���{��xg�����Օ$Ag�|����Rfo$��AKr��7�qR�lmm����@=��-�`m���?��#Og?q-���d2ߨԖ�p{bu<͈yyd��������mJ�������׺lzi<@I����B��SS���BK�K���Di}9���VH�������	�W��؃�Q��`�%sai�����=xܳ+v�T�
�L��b��ل簐��E���|���,��X���@��j�N%�4����t���sթ�;�'�n汯UԨP)1���h-��}<���{]N���qn������2����K���~-�����f���egV�W��$Y=Җ�������\��� �(�����Dt�ي�=����Ys�!�	�����,��Ũ S,Nu�6�h�>�B���)-y|���{e�FG_��JF���G'i�Ěy��ԌU�����k��3Yu_�J{�;C�&�t��C�';pPF��B������h�i�ō��y~m��#��=���ڑ3�$�W�وP#σd��|�e��Cՙ��Kk���t��]NO��d���d8���p=�J�$�ϵne�}��]m��6jN���}��l~MY�=�Q���P���˼���E}aǓ2!:��O�s��ͻ��ʠj�@&�+�~(����9��Kd�
Y�$�F�Q69QBJ�'=B>���q2ac�Y��)s��}|��!��>'��O��"L�ê��[�c�G�m���S���3��Ůk,���T&�4� �gÄQWxz}��l6�׼�����h�^(d��(�h���W�l��裻2;$#��g�@
��c	���N����9�*�l�� ��)�{�:���p�O�I#�t�����,,C���<@�����g�W\��A�)?�|I�2op���k k���Բ|�T�M��|Mx��"}�=̈(�2�aW�x�������+��8�o��s�!N�5�|��(.�����5����n���m�Xc�\�pHOK�f=�s��cNn���{�u		��J�n�-,MuA���|#q��'I�c�(#�K�/���z&���ߪ/2GԎ����Ĉ�n��I���J�vG]?�d.!H8�c�lhoo�����I'�� �^�#��1���i/��m`�kYj��	��p�&yg!!��Xb�~��}2��{_ǡ+�{�r���p��W�n���FP-?jF���Ĝ� �]~ɨ�;̓u	]{ak�B�߱},�z�>��������edn�`&"������ U�EG�qb�_
�9GJ�#��s=e�F��ÊN�j�W4����б�5�#Vr" �7#0Q�k����w���l����цh���cc��lO[Ϛ,�5�z947Ɣ����V�K����0��ʳ��"*o����ܠC���/��[���
�1;��=�i"�u|rCs�1<<L{9����HC}�0��E�Tv?.�$�?Oy�o3�+n�[����ț�i{�m2 n��Y7����p�㛜 �z~#��3gc�)��餤��9&�z��t�:ZR�V����G�3�]��;:SN�R`��^t��������s�	�Y]�)-�nnnD�C!��:�113S`�5:|OWUU�;ƞ���)�0�I&Ӵ��"�~�g��d�bPm4�0|<.�]c�C�CS}=ǘЇ�w��ȓ!�3�[9a+��ؓ/X|����=���6���$������s��M--#�x'QCta7��O�K���ΑkS��ODD.^�(S���2��8�НoH���*}�>�3�X4�	��kϠ<��J��h���+�<�Y�[o�d��'A�Ae^���8住��mt������n����)r ��D36��CXJ�%�ȹ���M(L�`: �OJ���~�?{m�gOc#��//,.�g<R�L���Z�^��j���'�cA��m������Ջ��P___��56(�(vW�xNU��١�͖�sS���F(�.wO�'�B����7����3�<�4$,3����OЍ���i���� �����fV�r�f�9�5%���2�A��T�&Y-�e�h�ވ�r?wb���F;b
�޿Ő���BMt���=�qYY�х�i�*@ƥ�N��Qn~��큨P��Z��ˢ���qRҘI
��G�_ �##�c���7���W`���4��W�$�x��#���f|n��˪�J8]��h���J�v�(C|^�ڶ��jг�y�����B�d��v��
G�N�T��}��ζ[I5Rz�]z/�n����
 �s�c����}4�������d��g��-�A���������rv��U�;
Տ��A��9�����[Ǻ��}�k�%�����x�5v��7�ᚐ��A�����+&����L�<JByͣ�@����C��	j��眢�0�#~l���#�z ����)�����n1q[��H��E���u|r��c��Vp����G"�+q׷�k��:(��A6,Tkn�ύ�Z�mx�����ш4�H'rHt�����9�@��f2֞_��t`��nw�ˁ)� )�LL���mo׈HH�������N�k��?Yq4�۸������(B|�n)O�iJ�vqBE�>̽Ш [9p��4xA��r�횕 �C�&��O`�����N�5��H1�w] ]ݝg�Atf򵏵��b�x-r�c��vŽ�N ɁG�`�; 
$yDhހ9�)	���7�|:h�����r���k�=E�]�QR
Z ��S�o���Y7���Fq�ģ厓��X��*���Z�is�;;���@lR
X�\[��﯊H�I�y%}d>�Ň��{�sOr������3COOLJ°���T��`<�+譣\w�q>EO��L^���G�g��㣢���3��!D3��&�l�/N�q3��=��*�6�47����?��{�Y�Q�ڔ����|PÇqt��N��@�5uu�wl��d>}Y>P�v�9CV	�D~�y8��̰~��8���/�99�	e��t}��w�#�D/q!1h~���3Bo��$�P�Hlll��M��}� 2P�1����m�(�gGF]ݾ#~ثAV�u��Vrŏ?�||�v �%��oT�Gm���߮:tHoq��p��8��b�����uu}�4��YH���u�d�+j�>;k��`*3N�Ԗ���uX.�3�\&*1�#�x����x:�n�������|���9cV	�1vB=�J�8TL�b ���3�A�@�ڽ���-�WA�� Y���wo�J��˨]���_�l�TR�]�h�			�D��my�s��$*�X�rНp��L�3V:-�l��2(��_��*���q���رN�x��P#DD��\	�>]�~�A�����-�lH2���+@ѝ�w陵�[��oe+����7FV��|�1ð����]x8�9�A�%����x�}��0�iq������0����9�P�����ysG�t�ɓ]5z�V�}��QL��
`�g�/j����Ȕu!��y���I)Ǐ�C}�XX�V�Ft�|�ʩ��C�Cz���"L}.���f/�������3V���թ�W#�m������J��b�s�D1�m(	��K�R�� �	��3�,�q�cc���F��hkBy�?��� �ş�y\f������w�sǓs�?FlHA՞	�z7N5B��N�R�C�$�rJ?b� ު=)�nrz�Z':c�Z�gW����J�\�.--=)��[9��J/w��w���(��#�X�i�_~GP�+!����X].�����Ж�'{ж���5��-�Kk���[�kZL�p�:�N}&ˎ�ˮO:��+�<�EFJZ���Q����S�*�	�.�%RT_�*�I�}��!w�ڣ�E�lu1�0I��4��c�DC�JX�Hu �2�SˠR]h7HA�����ͻ���|��c��O޺��q��-%qb��O��JG��҉E�ռ��X�����k8���^�#{+&�Į�� ����J� -�ڮ�̟?s�C1�5@��������y��
�K�Haa�z�J��k��:�{�٢��^(5
Vx�����fӄg�����)�c	1�>1Z�Oع��@��М��\BWƂN�:�ݑ����t�ܹ:�gJ����9 ¿�������r�(�u�s�=���Fe5:.Q=2�KI@����R˫�|XC{GGC��旕��tGWz(�u�<��(<��b`�'0���RP��sG���C6X��g��S��H��9�_���NH��N����L�WP���q����OM�Ał1�P��!]�9]V�2�+�u5�G"�\T���(J�U���妉KbVl/��h�v�Kv	?i��/"Ym�*�]%��N
��!�0*��L�lD�UbT<�������'�QS"�����-6rs������WD�Ń�cM	�_ �PbO��0#C���^O�b�6��ţ��^�xFO�3����N-�Qn=�in��$*z����ĉ���/3h+!X�|=�$�sdW��8�/���_��D����z-��P���Ꚙ�f�����@0��4=��'7����~��Hj�F��R�A�������ht�V�(E��X|�G����m4ᮭ��3񮯗�n� ~1t�U4�koL�#�mV�6\pvmJ�?S�~��eٓ��Q@A�U_�F��A��_�d#)�Z��k��p��=�4�1 �9|���F������+xy�̶`34��zD�&_�~�]ܯ��|%t��NJ8?�C�|�E%F�v�-0 ��S=�4!�AA�V��C���l���abFX��\�^yCT�u�ۻu ���c!~��������|��mj�|�C�m��-��=˴��d}��֎<+��0D��]Kj���2�B9-����G�D1Y-�����իW��|Gِ�P������Ru|�z�H:�rZ(V��nQ�¨�� �¥��yVr@PZ�-�c�Kݏj�O�_,�q|�G�Ca���r�/��@I*���]��6+��F���L�5B|�K�[����5���Ͱ�y��4��j�`���W3�ޯF��y���y�/num��)<���ϯ~���	wu�򁭔����Dd`+@�o�.܀���`I[�޲�5R+��Ԧ9�*gm��P�����X�>��Q��W�T�%��A�9*�v�A���Qů_e��y(�+a3��X/����?�r�I��*I�����0���;��e��+������K�%y�n�w�ܓ�=��S��wLLL��6�+%7B���jv�4�4_�1v���2�Iq�C�(�ت՞e��h�SN((�(����:nN�I��0�0i�
Hj�G�Z��h������Fm�pJ``���Sg;2�����7_ؾߑ�2�ٖ7B�#sz[��`���'����(�ee��ra�º��� ���G���-)ö��-�Jc�~ �ՅǤ��k �[��sef�2+��6s�<ljj�v�N�1�c�[~�M����dy�%+�`���/	��4��z�iM�V,��q��ͮ��~��U>O�5C��V�m|���|����=�?��19�s�ZrTRP��Sޜ���N�6��T�z=e�x��F���|�/
�(	����~R�Ь�g���:<��F��wxTwJS�����ש���$�n+�(~���ӍP?�c��&�Bi�����-��#�	����<Ǡ�趝Fr(b7@S�s��T�N���QV��J�6�&�(���d3�b����d���\}�S(R����9ȜR�O	�5�[ݘvLinV�qœԲ�Qw5�C�լ��(|���& �M�9 1`�������ث@%�v���؇7��7�g���.��;�U���cĜ%pC�]�'ʽ�b'644�ՍZb@�����4�g4�#ٙ�W�t�>A���^����w�%�?�Z�շnbK�N����HK�dy�Z��������Eս��cAq�
�}K�;+vB.Ǻ��������!렞�Ki	)�UA��²ZB��FVhE4N���@�9�ҟ��\ʲ�F�qQ�STT(���S���t�+W	ԯL����.%|0������ORQ5����#u%u/��+ U``22�����_�����xG�rJ-I�#�g����������8B�Io��@���.�����EGІ�����8hN�z������N�<�]��� /�k�(�#o�~)_���#q4Y�k��#J{|C ��m��K����h�
=��z��� @ę���ܺ��z�GbV�m͕*%d�i����|{{�|�����h)l���'T��m�lB蕇
;j�������]��)�ո߉C�x���ʞ��6�H�h�:��f�4��v�և.T��ӓr��7__6E�٦@b�T�ʣ�mŗz			C����$��h7Oܛ
"��a��Q��+t�b�;_5��˖q`R�����˰R��u�����d�\���s|������\����������O��Dh|ʴ+d���Q�OJ����+��29è+���q�?��9�L�`yf`lr��q��%=r?za���F�����f@@ P�C�g�N�M)�K�����/E�x�k`F��䌇��,��4 bk�p��ݛ�S��#*�v|	��b�����j�ƛ�T>�{N�D=�d�7���ߤvX�V�r"Uy�	Z�ǜ�$'�����ӥ3��J����c�XI���k6ڠ!$��z��Ot*�>;.���`��3�̄�@�C:����@�t)Z�^���
���'���!��q�U"E,�I��� Hх-��|�v��]4����\_�����|'vj���6s�פ'�R�-_RR���4�����`>�~�?�4�]�v���x`��."/	��	��� @��"R>�� ����F�Q_�f�FuЅ��qڿ�Y�#����w�F -���&�9II���鹌�����$��xy��̊�̀'��]�?Sz�L֧���LV���ɳ�Om���Lsr-AI�N��Q>P(�e؞~-�KL��)��T��pA�)�4X`��[R�@
A	��–��OQG'6!1Q�0ܤ쎝�_҇���JJJ�z=hioOpvv6��"wNHH �w+�l��@C�C:�Nww����RHq9�,�q_c]�^ZK����0��q6����4�O�Z֛��Km���B���G�'ڜ� ����/w��5��$&$�fs��:�2�UH��'�n�B5S����QuM͈m�C��"l*�n����M�ލx��ɢW�WI���<����Wkn��;8��u�ڃ=;>�:}�@ثءm�H��ڔ����sz��r%�@�R� �B���C�bo�U�d����K��N&%|~KNu�L �:l��<����c�_f��䱛�;̔�RPW�W�V7�>�_H�M�^Bv�2�s(�PO���܏SN*�,�ߋXv[���T�?�g�_A�y78NEE��۷7  .^���Õ��N��;�N��.l�:�1Z,�aʃYIPŀ6��5���B~oSR.HW�?011�D鞦�Ǥ	pi'�+������gY_"�5�Rd���䃨����Ea���G|*eRB��X���B�(�Z�M��`�_G���D��=x��L��	9��6P���^%ˤo�᳄-/�!r��Tt�� 64Y-;
ʱ��06m�A���}�e	v��1i5��ߢ������`�b�'b�;�c�9 x(�����t���!�<� 8�v�ѡ0D� ��Ы��$"�k�_2���>;T=����w'�*�i��1y��l�ϡ�������74��#c���J�;���:0֔8 �5�9e8DO���'��ْ�a�\:t���7�C�|��R�/�@e$�<q�壘��}UZ]V����"WL_�]P���..g��
5uttZ�~Z���Flfs�7��E^E��2���/Cf�OK�/-��~��;Z��q�5d��;j9EE�����~���_%���A%
L�d*!k\��U�{J>VS�J���jEb>v��3���j��0EԎ܌�����pVf
��*���Y��ݩ�<�߾}[ Q�*2N�*�Y���uy�k�5@� a�J� �H���&/[8�����/[O����aWQ.(Z��Q�?�Y�%��h[�r���oz��h��'#���"$�����UODzmģ������,m���B�/��|�D��|��Ѝ�b��/7s�ߧ
~)o��H�t�{��@XĜ���T����4�໨(ZTa�|ka�bi���zrϞ=��FA�2����L��L��4�F��1�r,ʯ2�������>��蜝��Mpp��Q\D�'�Y��k�8�M�Aك`�0>��F�egy�=�0A[EWQ�C���Wa��~��c|a�˲'��CO"P��������{��	���(O�C�y���߉���=������P9���M�T?RRA b�3�YA�>BC����T}���0�4gi��LEz�J�|"��LWW��S��UEw��*�o�9�'e޺}�'R������c�B=yx�Sߏg^��
`�s2C�jc�h3�L�+b���Z�L��Κ�!�	��T����������B__������:R��"+�ݷ�1��y:��31� �@l�HM��������w���?7y����4��Nԕ���,�n/�J.))�)ݠ���NI)aӫ���x��v�5���]�e�3�SU,���}h{�����z�y�������1�A�A���} ���WVVFg��1j���X��`?��u$a���:�ہ7cIv�3M.�6H�x��'0�Q|�yF��U�4D�E���`	����i�����<�Gю;����V���(��9�`�P.�����ee��b�-�ey�c�A���8�3
\:66��`�5�G�X��|l���Z�+� Ғ7�iF����������I(�A�>�rNj�@(����u��R�$�]haQ8�k�-~*�0@%�V��vL��h	x�X~���KJ������8^�����Bj�=�[��~k�����^�Co��"_]�@t6����4���՗��)�W�K5���fc�`f�h�Л�ٵ�LR�4�ڛ����3C�w�x�@ر�x�X�L;rV��+� zM�T��'w��˗��9���t�jI9�]z��X#j�(�O��������=L;~r�]�Ә�e��)%��v=�Rx8U�#㸞=��d�@� Rb���^w���%�͏��g3;�p�#c.�-%��(l�Þ<م��+���-��p��O�K�S��$��Đ�Gl���ag'�u �����\O�^D?~�3���C�^��y�������춝��	{�'A��qff�׊���&�ik䋼)qV6��M�������.���`逷�"��\ꄯ��羧!��K3��e g��O{�cW���߬� ua�ʁ�PiA�����v����7X����*:�B��J��yYL3���3��u%Cm���ϥ��W��������:ᗢ~C[�Dr�Ŕ	���iء��,��a�V��z��u���P�s�)�,�P���"�8�.��Ѱlm�0E��c{-����y�g���N�$&��OOK�^{����ma-%�|�ܾ�{��P�M%�`%�2=''��R��E��'���
���F5�Qt�D`���[*r(}G�5�9�%板���,9Q��������P����HQw�4��X��iӢ촐�)�Hd�6��:���D�۠���"[�d�B���`"&M�n���}�������������s]���y�s�s�攚�e �'Nq]�ͳOJJ,�`0V��8�&M��S��wϟyׅA�B���{�H4��}:t2q�5�uu����7﹤�s{��Ś]e�{��~��܋������.�^C�O�ޅ�}���C��?��ߋ�'f��+ݜ�?��
h_�\|��|���,,j�[<�t��F�o��׿���O�P�I�	���
^��OwA�t����"�|V��{xb��i��N��
.�9��]�>~|�}L��-�!g�B�|	����q�����Skk��}�i�������;oL�>D��fU�c���p���"_±g��f��K ֑����޼A���B�I7��ߵy�1���M+�x���s}vh�2��]'!q�̻�|�}JJ�ϟ�rL�o�_
��=��s#Ӳ$��>��$�Dz��mI��p���m�>�:pP��?���.[������~����As�i��+T�Y#`�Ho#�j���/��W�������kfM�Bs4š:7$a�����#ϓΟ���7�Zh�e��?��4Ȩ��>ɱU�
%W�pGY?wh=��WY1̞ff�V\=p:n�=ڱ�н����Id�y��|�zB�L{��$�[/2�t�t��+t�<k��u��eK����A N7{ʰ�) ��`�̥�{+%))��ҩ]]���/aKu��~p���W�*WC��(*)1��={�2-��q��2?��{�n�)�$y�bR��6�h|_�숊>�A,+�mdl�g�Rǩ�b���@��'O>��B���3#�%�����R�"dn���mϐZ$�<L�T���7)�j��><�+�ܵ�ӻH��?ʴ��j��z�/����4$D�	���v�+5ㆇ�;���_U^��ڟ]�A&_��
��gӿC��3����rh
,��>Ϸo�f2�6*NxoLE��Fv�@�8S��,6�[��NU�d�+*5�T�6��Ǿ���쮧�ѩS�������o><��)t/����B�f��-cx��e]OoI9��9��Xwp~��	_M�I�n�);,�<�����3��NΛ(pd���i#�(U5����l/u�cf�)�Axe��Nq�[Y�	���#k(�V�v��\V��ٴ�Pߡi�aYl�b��;3�ЪȕKh��u3�\M��E���χةCZ�_�~���ϒ�`i��/ڢ�t�!eI�?P&���%��̓dOC��n��O�d�]�Ç��� ��T�sI롛7o�}?jQ�~4�<�[�y�҉�CO�6�z�z���Q��FC�����>��=�~�a�;���^g��]�S�~vV�Bt��|�QĆӑ;7[��9�b7�����1�Q�#�I�9g��]��5��ĉ�p����7G�bb�_�Pܱٽ5�3��rc:;{W7c~ݶpv΂B�^ZZ�"��k�Ii�%T?;5�R೑��"�FU���z&;�����bˬb�Yo��>>E69�Vo7���M]BB�_�屚~���y�l(�� sG������%��]���}������\�Bh����EP��rAn�~����""��3-B*m����@dN�U�g��q���P�\h�oim���˽&���T�.�ϖ�H���[�O�Q�ir�h������p�����:��A���R��` 2PRp��682�ao��~����<�ݏ{�5�䷛4��A/�;*�Y���,_��6�/�,dMZt�O�c:����ʭ

L�K�i�:�'���,b����&�S�E>EE�i�Qs�_�L5`�״>2���l���_{��;�TAT��l:u��w���@�uu����N��P����_8|�S�����2�x&���
ܦF�F��]ȍ���H��]_�7�Ե���,R F|懶b��{��rЇ!{��~Gh󈩮����C��_mf���W��|F�<c�~]s����h�p?�W���O��N�������eq���b��5��zǻ��(6����%�$^Y��е�W�F̍Wm^�����q"�H ht���F��X�����U:hB{g<��|{i�z��fDZ�Hy��f��l�r���,���F\O��0vY��/�S3(o�\��\&y�.�Vj��Ϸ��ii���L����/��c��Ɩ��VDPh��
C�Y�l+P��I����ݲf�(��{�U;�<fD����ŴިrZQf�s+t���^=�l�*պ�T|�DMU��Z�,˰n׵�þ}Pୠ��n_=�d�\	}bD�e����I�[x�p�z4[-#--�0S�ٽ�5����3VV�oֻ��m,��,+K�����Wf�9�����g{�f��x� MK���5UUC��^~F�Ӄ�� �4{T��8�� {j���.���_�=���Вl
}u�e�ʯ�,4ڱ�MKK�6��v�J(�˄���p�no�b]ج6����:h55�YU.t��7*kMo��j�x���ܡ(�Lh��jv�N�b�����}zb5�C��>."x]�͒�\�&kkk���y�ed���S0�,g�%�r'ؖ�,��N�N fF���>"~uX�5�kѽf+��Bn�,��5������Jq�,�jr5E:)ŮP9'?���PLD_�Sl�-��J𝬌����nK�,>��ْg?�|��e�������عxv�9�b�%�J�b�@�����0Z�QɅt)-O)�FZ~A�q��MI�������ʗn�]k$����H��;vUGmDS��T��Yi[��"��]�ot�1���Q���*�r�q��Z��\�M=$�g�t[ǌE�agl�����b��������kb�f��+bD�˽���f�ie�EE>+ŇA�Q,U��%[B�|�z��@�������d�-ǾK�p6�[���T��9�|2�on|E�g2)�8�R_���u���!_�[Wӽ�fʍ���WS+$f5���ʻ{� [��	��5��J��+�/;X��~��xz�}�kj*�f�N�H:�;�:�	Z�\�<��=3���/xU�d>�8\O�,�B>э|���0y��jϚe��1���*��N�)0�I t�|%,}��&#s!���T�GQ/�Q����;���\��\,B��ٯ�d8�m6����3�����
~$�W�i���O"	2�c}�g˂��G�$��q����X4�-�l�<�%��|���EƖ�k� 8���_�~��RN����C>m<�B��o����Lb��*9ш�ٝT��	�q�Q���J��ጮ��ж��dߥL%�� ~ii	����\.�=;���?x�(�{�2�������l�x'�`1�Fŗ�f��ƤYE���m����h�tS�K!�tg���#�:��^�,n�����D��v���P�A�
��K=,h�ۀǭ+p�Ӑ�aI��*u�~�q#�G�N�퓏J���jEW;^�M�Hr�K��s{n�J�dv<�R�,:~����s��z��I5���t�.��~��r�
�x0OOŔ�ҋ�L�V�'���dY؟��R�/��������1e���W ?�Ft~5^�����v��Xx3�6�5V 50%��(Χ�꓇$���F5�'��c���%�@�\��G�bl���[�4��8n�9`��jP�El-���p} J����j.�}�����lΪ��S�!�E^2�\Mq�Ʋ0�7+mС����X�%PʺDhU].���ͭ.�gǜ9���-����557w!sg$h����yЕ�뾮9�*fb��.V�&��Kw�6[i���%���Kmħ�B%�vf�3)I�]���~�7��/��+�*/Gr����es���y!��?��;�J�d�y���>ȇ7a��V�BB��+/����S�V�#�}|�fg�9��TYI;i h�D���>,���?n�.yQP ���~aC��_����&�=R��|��*Ò����]J��Gd���L�Vȣ?��.=��}���6��b��w����n���g��تTFC����ujB"K/�i�����G����P{ׯ_?8�hP��^]�^s�Y��?�oH���5�-X�WүX4�h�#���J4�E{����|tl�U5�͐宋Xh��=D��s�F�^rL��l�3 ��PW�+���׋Iayyy�H.�t�X:>P.�Քa6ؠ+�᥼F4L�,�$Z4�Z#�������[�+>{����]�����1j#_XE�)t���G{�#���^���h�2�����^�\
+r�5��?�#:�#4C �h����\yb5�)�zlտ8Ut�T���%��d7Yn4�4�mq��0�볱T	7o��g������3���"��B>�
��j�g�}`;�p'��H�w�����ć��}�QQO� �S�q�p��vW�@˓C��������U>�`^�P�V�!�1�"�*K$ދXB���A|�v�`���^���]Ǭ&q�J��s�����ٹ�����Om9
�.��<�@���=��h ���jAo�[�ԋ����W����ע��T��Ϙ�o�OGhXX�������,'7Wᠹ����\`��3/�1I췟^PRR"��p� �*�F;0vq�7�GD��fc��n�L�`Y����Q� `
�T��>��A#����xQ��DXU�� 
����͍�q@���@p=8��%뢲ɝ��MsS���b9�-AJ"]?kd#>�"����ѝ�j�Z��?ӳހ��YKۅa:`��г"��{����Jk�f�f��q���R���nk��6y,�~��c�xj#Mt`�f�ޏ1<*d���K��C��g�I�h��<�t�P�������U$��ua��0��Te����:��_�ܒ ��ljߜٝX��>V��Z�(Z�X�y�����_�����~vQ�˗������L�JOL��Ҡ�qFd@�C�݆��|�6/o�h�����Mv��l��1�p�
�1�I��6Z�VD�B̵�םxX����DT�f|��I#��r�@�^��y�3r+yK��XA���Nsb&S�2��4,�]A�1B�'�Cۡ�ܮ�213Cڤ�wڋE�pV��ݬ��E���-5�o���9o�9Ya��*��TV�Żv���B���$�pz_��4÷[�+��f���8ͭ�2=�t�����y��g�M���Mn88��.Ls�
�����eB��k����&-���>����,�Zjg��9��!���,��C�`���i����{A���\5%�[�TF`1�CuXk?�/ x]���J���U�9d��f���]=���Í��a���"��-!28��`g�#�0����&g���W��NߛϷ�"�e��&�J���ţMfHJg�N^F>�>b������/���N�!%���uˤ�����[�s�w�::�`���D (!=��v��:&OC��X#�g �E��}}�(�o�'l}D4�j�RW���C�M!��jܐ*��35/��zB�[�T6Q�&����F	T<3����q�=�L��*{�2z!k`�989	ZrB��Sj�c��M��U�[w�M~q�����:��+{R� �Z)c톱�A B�X��Ǥξ��p����xvH��G.��������:}��ę�2��*d�֗�ȤN����W�a�aF}U3pj��_82�Z���-!03��0�e��J�f�;ھ4�I��J&Rg�.N�|�~SI>�	����c���s��A�7�{���ПiQ�Y��0N���|Z1p4�����^�fBZ��6��hbzbx�z[V��܋ə�V�?cR7"���/�rB�taf�ƭUFFF����+C������w58��a!�_��/��N����RȖ�. ӻ���|����A �Ρ����&R�nZ��[�!\�	�eMDx��C������H��E�E1������g�0$�8a�W	��/�]��:�C��k���3NE����xa�Կ�|{W�R�m�߽2,+���(���Č��0:������j��eB�X!� -(_�!��v낏}[����aA:�z.���WW�Rg�R;�H|��ya�o��U���+r�V`o�a��MC���^��V�
YD�b[�ཙ�AY�X�di`Z�͞��������{ȣh���w B�r@�Fŵ1\�O���� G�K$��K|��?��t��X�h����	u(�`�!�Pc�w)Y���s�D�	2���$5��a%>J�VeRHW���G!H�YQo{L�B�R.�g����Ճ���7ЖO��KCw��-�ҡ(��OS��@ 1.ž�R�1&!��)o,�Τ6R��<iYV{	��m�1�@}�H����{��v���T^��:�P�����U�[���@k�Zc��V��<&�_����$7l��p�gU:��a�*�Z��PA���_�DLf��Zo~����{�0� mq5�*[ qM�Kwu��,�������[c��$D�󽁢ET�2-��0&5��}�E�%�l�	�P��b���،��z��h���ҳ϶�C��YM���#B���~uXmd�=�%P�I1,X��|��Xy�"�7�2����BVA#7�i���ۅ�n���?2�
�&6�6I��T���R��s[�?�
���T���Ŵow���J�����Y8v��p!�֗�{:�Y~&��5�6��06�V��}�-��+�I���Q�������s��;N\zCsy��d���߭=�oρ�����!�ϙ���QV'���6{&��c���㥁 ��݉��"U��\j����ˣ�!&n�`��oe�@˽?N�a�I�/QD'�@A�s/�Eh0O��{8,�t�������T
����j/4xX�i0�=�)��;��mr>LZ@xK�ݡ�`5ǃ�B��<U� g�󓰻�84� W�B֝���s�%O��s��w"��{��r���!���>�i{y��V�!��W�F��a�L>�>MK&^؈n���zM��~T�ݣ� �Zh�a�9��=�T�]$<#��\�{�RJE�����!��P>����U�9��$.�F����c�md�Tll=�AQ���zx1�a*��'�>�<#U�<�����r��{�zH�J��>B�~�p�/�"���r���������@��w�W��pؗ���o}Rԃ}�6���8��IdxσyZ��|�����_�kYs}O��Q߁�ۭ���)�~3��H�/XB�v�.V���{>{o#��#%z�סd�`������6����?3��BJJ4\��O줔#�X�I�=�@	�6A���Y(�����7��ӚJZR%�)iis��^�!����S�*PwU6���x>�})V����|1��rix�9���z��(J����-�0W��b!c�R��J3<����3 psMo�#4�t �۞d��m�Sf!��XAyP�����<G=�B|!���E��_Le�6�=Fhm��������e��E����=��{y��c��������Qb�o��掦�cr8��|��Gx	٫j�2������V�Q8��rU��w�W�(-�/���E���=�@0��^AE�@��(�e�0����¨	0;�7o��0<\�� U0��\��5�!(���N���-�����PT�E�=�B|�*�Y��Y_�������h_�J�Gf2m���u�x'8 �l&.�
�V.�ɧ���\�)^ (-�ּ�������F���^Ed����O}��V3*:����w�"��l������\uW]U �	/,1� �S�Q]��b	x��M���R>h���9�KvWk��U@c����ۄ�y���Mqɓ���ˈ~L^TT4ΑO��[���-�ar���PQ�	@dlT�@�KE���fm�3|	i������x���T���;)�V�@�WP �a�H��!j�P����"���e9�Y��ɿ�e��JONK�G��j�Q��3[Ξ����z���� ��/Bh�&�"'�*6�e_[Ȣޅbƀf�r��O4{ ����ٖ�j�s�Wj�mZ`$a�G������$��p��#ڮ5��oϤ���$���&�s1m
�q�]�O�.��� ��ٳʿ��\��g�� ǯ���^���\�9P��X4�,�$��[N��E3 ���V��!\�Ҷ��*&uˢ�?w�4�A��,ּ����ݖO}�1ߑ��+,؀�|��͚����u��r`T����OV
.  ���Ѫ�u���\��o���|���^�#"U5ፗz8�H�(��g����,��^A,1jF���DZ<�<�0J�1	�7M\0���<V��ym{נ2ς�b��FF:sA��,)���,?��� �N��OӶB';�T[C�y,0�}[�&'���<��d�XHY��,��ZB�*(���+�7b6� u[��%r�6����~+wQ�d��f�ӷ��ʃ8,� �j�;78O'fK��, X�L�����C���?�E�nw~�"��#B}&�&?�0]C��d���']�q�1����V �^{Zw��Ql����z�w��B:��(
,������!����'�Bl�
��e1�<���,�£���ַp �``�^�푆%�=,t-��nf~��R���"�K��9`�[��%4�v"����D�	i��ُ m�K�����N��~!PP52�F�v���r�5�FǢ���E�
O�H�pl b��F����5�@�f!x 	�Y ���fH����	��* G@S�b�-(v�ᒁ{R�?5%DDm؈����A���&3��[P��%@�Q�I�%�� �,�.Q(_��w *	c��EA)�k�>��S]��⊢?E���o=���2U�nOJ�+��z{H'=m
Lbʍ�E�؞�y���7S�P�A�n׉��k�\�-!���P%�D���S�� &�"&���_'}<��]1�$}�*�Aޖ�pi%�t$�$�b���>�,d�qEO$7H_U; '�ٽ�{]��5�7��+܀~�O½p�Y�W�p�/�#,m��Y++_�'4s�@����s��Cք��!F��KKS��޵F��S:�
������G�7��"�S���eEb��PD�Vpm�Ij��,�Zw�.��u?E�,�/E�d2g����L��-7�n���P�b'b�)�"pX��"�け�Ra[�̶�Gܼ��{۞� ��'��hP�ٓ|Gί��c�Sߦ�w!�n���5�/��f:�4�V/��#�٫!��]�?ձZ�['���� <��+�*K�K4��BJ�QQtfvfi��~Q�?���n�1�̜y��F�޸�&0~j���5%�.tp��`N:\Pvl��%��Np�U�r�".���%�R�1����Z�U,a��7m�_�����L��ۨ��̊>F��h�hK�OS@�UH�N��N�8��Gf5Qг�tY�&�I(ݳ��xm@����������Npf����t�6o(ż�PX̿)�Ǣ�|/A�@�����B��hy�'�7���_L���"�� ��D<�w���͎�>�`n�%�Z���p��}����uut,Ü<|�Ù�!zT6Z��Ӛ�XD��"F��Q�FA����B�=p�^��=�@�NN�ߗL����:��m��<��psԹ��;�v����0���;[�k��;��)of��H
oN���1@��3�<+����<�n�o �<��3�tͳ+n�����)����4������?h�ߔ�M��Ԕ���vi��49�����bn��N������:�<������m7%Ο������o��/M)�·��*50��p0�^c��^>
W}��{�C�����Х�.d�����"99٫jO)'xw{~����}������1��C?�#�,^~�<����	~�GUph��ck���ח.]o�̓�:5�}!��G��%���em�GS�SN���ܜ0V��Y��gZ(��gu$�T4�M��%>���]��9.��GA�}�h���v坾��YB{�v��W�B��c�������~cᨁrҡ�16�-���'�,��1��6MZ��{<������ڼ�Q�?���>ބ��?�3(�稷��N���x#������`�k�k�����8H���U393k��D�XL{���;t!�2��6��x�3��G�Y�͛����Д�n��w�4��O�%n3��J��|*�u��v�C��L�4y�}R�w�(�K���\��-�wԋ�&��tV6������Ŵ�OI2|1yO$A�|S}��7a1�x�W��,���Q�&�חx>#�
[�O�7a����.��df�I	�����͙S.ڟ��2��{2��X�ЩX?/���Us�J��bӝx"��?_�7����� O:�t�k�E�����|�}�R�D�~
�S���?
���(XL֋vށ]��~��%�����ze��N���3�C˿<DN�^~n�m"�u�o���2���ny������kGd��y��Ky7��?�J�����?���g��_<=�kk��ԄD8� �>�SQ�	?��E��uM#�\��}�� J������)����wZ�o��ۏK
��x����8r��Lv9#�+_��ZB�]��PP�m�ޡ���D�c`�������Ңh�)w�ܒZиvA�a�$�?�%���.d�W&����ʫj	�bX�y���ff�@�V#�$�X�eBƲ���Ft�T��1���NyJ�*%�N�>I����E0�^,&�}��?z�iwKEpt��� �q�l�3?<<�vtr*��= 0^�q	B��u����o�����.���r>����q7���,������7u,ڌO5������Q��c��/�P[�A���Q�d��HUB�?���t���*A������L]~;��wh�h���x\��ܼ}֔V�8��t'�Wj_XU�$!K�e����%/3V �˯;&��A�ǧ�6a1
y|�v���ڻy�~����n��sU�b��_�M/�iiq��"}��7˿ՠ]��[�8�ay�̕�Q�1�/�H�t>���!�Qj�Ӛ���}@���os�ip����2�Y��������F��>�n�Y(�Ï�Vp^���`@`FYoT"W-衆�`�����i{���x��r4-��9ދ]�rO�l�-���s&�����du]zެ?���z1���a꧂�"��I���~�d��2^RT]�n6s���zM-Ai]��#5|lGq�����r�^� N�(���#��ި�H0˝={���wI{Dy�d���Ӽ��#ɶ��%��^-a���l�J� ������8,�J�Em�6�n�DM�4�t̜�n��>�P��:�5m�����D�KА!�B����u�)�}-���T~=~��U�ߠ$���_L!��S�5i�%P0*t��G��D*e%:��E㪷���_�y�߾ ��BZS��&�/������tQh	�J^SVYЉ�k
���x5���ua������'�wp�1� �Ŵ�Gɤ�����.gXٗ��!:w�Y�[q�xϾ�W"���K�a`�u`��`�,�
%~��ؔ�6��_��+��_�~�~n���]�z�,//�9gi�hևf���,ֿ;.F�[sY��{z���B�I;SS�� {{�g��%�Ѵȥ눃�c^��q����o!^8...��˯�B�β�����;��F3_[��zG��Ƿ�]�G�ߓ#x����g�PЫ�0��#2zz���A�6�� �\���55���f.[�
zC���Z�#��`p'��9��a�1y���I��yMj�J�i_���N�[�p�g�g�-d�Z'jiWD��Y���Lr�r�z�Z}Uͧ�4��o���΋Q�/zc�'&&:B���a�����(-�}ݛi�ҕL���V8���3��i݂��v=ƀ��n7Xv$K��̉ϱ�U0V�ēL��V�EeƟ#�SA�Nv��֨&��5������N�|��/5�i�kwuԶ���ZV_��6Ô5x/|!b�;�F|�A��^Y���S4%��gS�A~0ӺX�4���=p�pi�=���0�����e&� �TO���t !�Y��t��i��$�LVv�qb��G��G�î�=�C� �>�lr��������|�4�F[�,���5w��yjTXT�vw�yvW�R�R��6����e�wvc@����NiM�`ɐ7q��IȆƞ��23�h���ր�f�����gr-�g�AU�9�aG�c ���+���v@��h1�ѝ��3��U=��H�S���!C�X*�9���/�Lc�@Y�&�X�W���U���I�}��ZZZB�
_s/vuV�f0P(�섩AV}z�y~y| Xk��7�͵Y�CXd�*䁣�YH���=}�`�55�J�@���ҫS�~S��I���U��č�y�<i��1�i^�;�g�5�5T�83.f��6М8����hݳݛ��5X)�<����L�t��q>}8,Z��5�kbi�^�CM@�ib��K�&�cl�܆��0d"M���f��ԅ�����V����V�2�u��+a鹝Ú�D��� �	����>9�o^���5X��������N�5���D��ּ;���6�*ÜU��0%��u��.�hfV^��?�)Us�ҥK�>-P����|+QQ*n��7c	�u4D���0��Q��Ty��h��Ma���j�_y���Ȟ�9�����?�%��X��%�ld
u��>����ߍ"�~�7�!Xs��8U�']�>�>��q3N�=3Ů�ג՚�'�P=wl�^�����xX߼�{T�߀.B}�$/slj�,�4y/=�L���E]K+`�L�e@NϚ��Ԯܤ�g�2G��t!�D>�^6p5^�_���~�2:�3Ͱur�]i�JN��N!�>�<�L���oAB�����&Cw��Q�2tْ�SX8������L���ʛ�6,�'6�]��q�t;�^7X%p��u6ͭ���HSd��/��b��q�:gz9Z,�[��l��w��MK�6�H-!�H��1:��؆��I+WK����)-���z)/l-T��f�l^�vIc���� �,�
�;у�� �&{�)N���5Qtu#�¢����X2�N}�gw!{H*++�}�}�A�@V�'C�<`<����3�JʾX�b����2=>��
_��d��B��>}���S��ѬQ��Ǥ!{�K���N��k��֣< �=��ƐH#G����).�ye�I�[����KQ�~�6q��S̵TI�M�	�����~	`� ��C��_Z��<{���Y �];�^mМ�(�JK}����`�X�E�p����m<w`h�U}�G�܁��Ԥ�;����-=== `�$��6��s�������s��}@�3=n�'�~���uX*`z�{
���2Q �^G����(���$,�F6B�#Ѐ����.C��5�EY��M����&|�U�I��)h𩏣pӄ�]��W�����Eݟ��W8����?�O��F4���A��(Ih������(7�.�2��P#���PY����2�׳�>l��W��!�F�ͽ�(��3�	��k��¦E]�_�~��u���+}��1\l�t^m��ҷ�(�䬲�1V�>�ϵ���n?{z��C��p�V�����7�Q�r+0��r��3����a&�9�rZ�OB;�c_c��H��-%y�w��߷�~Oc��AF
E�P�`=L�ꃶ��"�څ�N�0�Y��{���[��������m����n/ŷ:�ܱb����ML~%�pp������(��[�˺��Rʍ^8�Xi��Q�5��C��%�%^C�I�j(�@�J�12�������(�}���!��-k�K���mɟ��-��W�@�I�hF4hf���
�.�TT�C=��$��Q�ԀV�k��F�R� �}S�
� ���m1�f���V�t_�$
/A��Ð��9�L�)��n���[��IHJ~�G�]�g�ÈW��S�)���^{�OЃ���P����")3c�`A�tK[��T��/L�ϩ��p�rBMM-OE�P��1�҂�YF�6m�<3��z`}�rXߚe4�rQ�V}9��9�s
_uv/��j���Hp��ڂ����gA��c�jΙ"�2Q��UfM�����AG��e;x�(Q�~��*�6AD�Km"�']�̍���6fU��P݄�1�sz�d��k�5��@���j��=�U�dV�摻vU%@EWCĈLi��h�?�	7����2��
�V��1=�Ll�ѯ��V�ڲg��j��TR2�c�4Zw�<^�PqK�ak��O��>��ҟ�ּ�
����u�����e
2�'�l�$�4�?�9Y$ؔ ��VVF�8�Y��o�}�Xt��l2B��Tq|*�G�/Ͼ����K��5ss����.�ӌC�D���@��t�*[	��hǾ�|g��!�$�O^������I��W �,�$U�$��/����r��O�}��f�|v�g����Q�@�(�G��u�-Wj�������}��h�k�Ǧ\��{�� UN@�;�tkS����^U�L���O����
�f�ZWf^$�?
ι�b�
'N�;��'�Al���.�q:=F���߃fc9�KTϹ0\��t�ji���|�@�q�ӂ���;��s��� A��ck)��a~'Tɓ�پ�>}"_�@��bS&������1lT��W���XL�:�$���e�X��d�j)L�ٱ��}ך��2�!ٹ�1cu+��'i<����<�T��~�����i��lG� i�ް(���/���`���R&r��08g$*Ůt�L��w���� � ^�p�e��c,8?c�ax>�Pk�|%�*�&7��؜Q[��9�'�>���v�'�]��sI�Af�[���Db;��B>�px�I
I�k��q 7NE���%}�˯@�(\a�c+��Sؚ.R�A��}�"�/
��'���}�h!�Ѷs{�\ў�����2��ln�Z`=����h��
tғ6�Zq�$W�%��h���7����Ӛ/��)�%��צ����dZ�~{}c8�p`�K�]l�L�+�����"��~=��u� ��i��t���â�r�p�l�j��t��V$��R�~<�*�Ni�����® fMߋ�����׭���K��T+���O��Zd'c��-�	�����n��3��JNf}��kOk����m�n��-hj��hv�JY1iȍ���� ����S��5���{/�9�N�
�D-Qa��T<�\��ZF;&!!q<����-"��Ϛ�XL�cz:�A����B*Z�ZC[������{���l��#dZu8�0�D$�m=��e����k#�T��M"R�p�!R
p�z@<+>�xӍ��I⿽�h�H�H�f,ӹ^���S�h&@3�N� ��k��ӕ�'�[�9�	����@]���S�<p��x��^�1�/��/��K
�ӽ��'�)K	��7Z^�ӻ?�Oo��P\ʕ��n�̶�ї�Fo���+��O�Q�,sb��<]d}4c���A�p"ǄO�p3Lw�k]��LO�Y ���ȩnu
Db�S�!�~$�;NUM������n�Ѥ��/�b3@�<~���mڨ�6_E v�H���N�2�^�k�؇�?� r�6�F_g��ޝ|d!�:�5��bGbG�?lA4F���1�����u��4o8-��
���L���	��EsI�c�t����`�=z�ś������ϻA&���L���-���l�!���Lgf�^��ͼG=�e���I9U2��M����:�,(�|Q���.�[�a�ID�'͎��r�$�W�/]���]��j��fS�u�E���P%Mz�9�������l�N�.�Y8�q�\��U5�����0�s��&��_�?�N��^��&� 0��IS�|�6�7{��]��Z�d�N��k?55UJLz�j�Q�3~���1,#���E|�i!�H۠³y�ORAȞ�V̳�߃�LQ���U'ARކڦ�����p��kEH�@�m����+�zj���ܾ7�(�G�+8�C����ҪFE��>ݛt1ݣ*��� �Q��'��i���deHr��@V-�ܱ��z�Z��2�ո����Ya��E����Wt�P2�Rj����.��|���h��eT��r�&c����X����i.""�%^��ޝ�ƛ�H�A{~�6�3�g
�z����A�G�m�9<'����h�����-��YK,p��P7!��� S��{� >$�[�=c�㉤�bQ�o���+�x��TV�`��d�����	��(�u���vq&���2�+��Ϻ�h&⪨�ʞ������
�tO7j�xq��>�쏄8����u�k���~nE̋�y������ q�������J�DYFW��f7���~��s躛ڳ/��S7�J ��F�z,�B��Y�R����B��"?��\�j#���{=h�ǻ�i���d�Z�Md��IY���f��=�e[eJ���O$�h�Z�����3������g��?�=��d򀊺�ff���K<f�*p�юաVέc�ЃZ��|�;��a����4���ܢ���20�̜�~vY������N���!7�<�Q7�8��};"qޞ��>>����t3pX�8�R{��4OQj7L��xT3z�_�8�g���s u�h;Cy
�[�m7^�{cl|��#����}x��S��VE��.��<���B.�}��Jl֩Hs�\��Ɋ *Ԩh��BeB\�,UaD0���-��DkY�B�����s�{��T`i�v�?n�D>"z�	�8A&}\
��Rl�1�B�.H��� ǘ�6n3zp�/u�E�X
�bE�4��>��~�J�
cX�1�䞟���b��:�',@��s�z��1}WMЭе�9*>�)�=7�	t�3Ʌx	0���K�c�*Z;�#���}�
؎}�2�VW&Ϙ.ӭ8۷!��]��Q9�B�T*+N	����qjp���83W��ّ ~ϓC�/�Kr.�7��!�O�w�R�d�dq����}����&ɥrxɲ�h�УQܕVH}E���T�eLגIj2�zP��������v��l���
CI��"|,L�M����Lf�%p���6�Dg �w��5��0kɟ� �.C��@� A��
��)qk֥��"�$����jg�@��#y��I:4���Y�Ā� *2�ھ�^��� _\H��� ���j��U5���
#�61����� ��M&iI�2$�w`���V�I-�J�� �LR�����%$�Q�I��޵�`����<���NB���ND�0Z���ǭ�	d��n@�֏��I�k�͞�t�kW�g���Xu��_����j0�b��:�F�����K�4�#���T���mܯ�<x����#���2�`Ц����?Ae]@�����\�}�o�S���!G����
� r�����]܂Ԩ;T	,��6m�B^spO	ZY�m�n�, }�f�}	�{�H�w����ߖ������!����D��f/i�Z��b���f��(��ϗG�H����VAB��ln���%�?���뵸����@�b���9ovJ�N��䑞n�	���Ϋ��T�$}���� �W���܋e٤!�XI�B�H���S��ЃM�q%9inE&_��\��uF|�^�?�����i�'_�nuvH�+Ю0��X�.TA�B'� Ө5��H�"�VTTd�^$x��vŰl�;#�S��I����Cq]��jB�U��k�q��f�! ��t��wO��T����a2��Sa�v�k95]�`&�5�Ї1<�p�⹫���+���]�&�G�����B����{x�k�L���c�-�.*����[�X�RzC�����V�Nh���yQVƁ a
��b��ќ�b(�IG�pX��;�b������e�q�"٥�1mRh�ź�����,���eJ��h���%
���}�,���vq.�����q��wR�B�J�h4�	�}Z�WO[��)�Ľ[�� r��T�`1�8
��[��P�!�ֳ:�N}q.��J�OԘ"���C�:��H&E�}dlL6�y�E���������/pj�L{��s]T�m@O��rE�+�e:�bf��!���<��4�8oSm_;m�2Л�Ye�'�L�-�}'`{c��S�wyYp#��*j�*&�j�/�!��9WLw�l�S�� �1,� ��
3��j�$�Ǿ�c�SQ��-@��i�n"��%�_j�(3�N����xiKX�J;���`L��!hOv2������m333
��Ѹ�� ��8o,��]�Ӎ��]0�ڿt+�]�&����|��zt+z�74����J���h�G��� }L=�I�I��޵&�l�9i+Y]1�^:d�RTxhX�� ��lgr�t�z�Q��� y�����T��c�Z`���d�"�b�C�E���u��
�'*���N�TD�Oa�Q��!�t��?�S?͢t���u��g�Z$�E��f�'�橡�G ��w�X*�,'_�����a��u�p���B�2����-�O$rI��s��(j��DL����J���9�CN�E=����)���{,�`���B��
���g=;���w���K_?A��3��t����d�弐L�~7[b����畗CH�N�¥J5�ȋ&U�&�\\�&L�Pe���҈$X����4����?D�vi��U�4���!�APA�%a��
���	�q��+�"� Р� � F�$�������eWM�TMM��?4���}��s�Kr�<��ƠM��'2���=W��!������ku�X;u9ߠ �o�5:i����Ѭܢ"�)cSj�9p\#�z��o9�e��,�ވ::4T�*�$�'�������_�LhV�+��97>42�f)	uq�����`������2hP
AE������ӵX�9�\�`�ms�O'�To����.��K`�.֭�ov�B�5z���:47�����m��|�CRe�"-�G�4=8%L|h� )*�D�ۡ�r�Rhe-�"��"݁�	�333�����_���^�Ű6+�F� X�"���O���D�Ͼ��~i09`M�c��c���n)���4p���6i�u���KR���T��y^3u�AcڍB܅��s������C��{?}RO��O�s�h���P�e�W�As;'�U��T�n��Ƴ��<H'�it�t�;���X�;��t����Gտ���S���-Po:�w��\����I�o@3�9�ϟ�=�j�-�8+�)ڦyS�]�-��|dg�
v~1��|i`F�mJ��Fe)g��}� �4�~���L�X��5��x��-����XJ`���d�jO���b���&-D3P��I"~L��g4�vd]��o�(��Y�� nL~��'H*�;�������|��ZO����SÐ��*�E��u ���~�߇�
� �J(f���޵1I#���i��4w	�[7�:�ʬ��r��Խf2�q�!z|p��+"�Aޡ��'��Z]]��5���I��^}ceip(�����6r$�W�Y��C���i98=����i��~��Pcj���	��"�����b]��&�q+��b�G�;I�`�H��9֎�*��Z�E�����!�<�B]_�W��S�066vy~��i�_�6V�?�fИ�Zo��gǳa����(~� �RHP�����t*�\��$�t5��ѸKpX0�)�?��]֜[	�3L����7��|9�µ���_052�5���B&h�'�M��}η�N�b�Wśf�1j�f �C���Q),�DK��@	��g���^���M���*Ć;)p���v�u���P�,�\�s��^@��|�������k����###��'4F���G����~�Ih���b�ξ��2���n86��k]�(����=�N��m�7XgD�2{�^�*��-��<�}�W?��UaO�}���4T����ƿ�`X� ���l����KGڵ���&>��X�`;;a��\qE]�_oc/�A*�ŀ[	G����9(]#��w�V2p'�qP�;�h_�]�n�>\)<\W1[%�yҮ�hX���^#��Δ���A�{�;��p�v�-���֚h:��.����!�;0�*뤣����S�r������j&���V�w�^�	܊�U���\��@�o����܄,� �9�/5U��uu��v&��ָY\�t����W�#�l�a��gw��ЖR޳� ��+���l�h,|�7<	�Z�x�~~��O���G �k�~ɣ��AX/FjdEc�;�[>K������[���4+HC@�P)��Z���!��Y���*;�	�tPRw���[�|�����m��v�1>�F"5��0C�_g��2S���-��rK�☽ٔ�rIP��ל���9M�R p�@�n�ؿW�f��{�bF���Z���~:8���xI^����[�M w����!�W'�!���O琤��Ҽ-�s�3��S��|�.���
��g�NR�|;8�� ZOD��.��[�Ei��P:�k��=&,EͿ����5��(T����`����T�POiI�ͥ:��L#���� D`�V�&�+qde��U�1t52*w���� �E/�(�DO>�m�U� ��nS�°���R�6I�nC(��w��e��ޭ��3K�`�b���������}�0l��_��������t�jw�?�!���}C~���t�Ƙb��K���4�Ǻ���/:�3���vCq��'�.��7��p���m��+W59-�>0��æ�ˉ�r^�ƫ��䃶����I�P�����0�Έg���������f��?��{��j:z�o�[�.�V�#���aNat�4V����J��4�n��c�rg�Vl�� ?%�[�=(^�IƜ4� Wq������I,����[ 
���y� a�I��	���b�z׭f���+�CK�C���y���X��@�DvV���d�q�~{�4B#]"yټ�d���6�5\~3^�Ix�Y"2��i�0��GK6S�l�n4��:�E��L@P��d֬_�҃A3>j(�����1�}��İ�� �, �Z�~X��w'���hc4���(�{���_�U����\3���n�+aN�p�.��f��N�L���!g���.��3�\�5U��A�����deА��T.��~���D���͌���^,�����XY��f�����%�/R (*j��FW�Fs���`�=������l����3(#%`(tC�G)��\��lx"v?N_�V�9GP�X){rk�dq^fT��d���X>�c ��'X�0�Þ����fH5��e�3�H_��cT���R��ߓÌx�:��8����V#�����Eu��~��,��`��@0���n��[�^���m&�*l��~y֪�pp�������L<~��_�P?
xw��*�@nb�� 5-+��	x�\wO�+��g,�Rb���	
**���C�~���(�2����5��"c;��*����	C�#������`��P�	)_�Ic-��b�?���ک�j�ik� ;k�6�@kn4����Ϗa�,1�cb�1,���c��MZs�ʧU�ޜP4!^���w�Lԥ���q�}�ꕒ�/�[��0gDA!�p"{E�?��N�s2)�Q#��ɾ�}[��s[��ꩆ��id2�5QZ��,�,�����N�Th	�p����T�$`�Z��fs�e�P.�4�ɫ~���@/��nU����ۉL�E�se�F���7I��`,_���z��Uׂ�Rv�ZYQs���=�K�˄V�~�L�;��̊�����'CmY�"_C��w̆˷��	'�Qo���F���_����+,*��Q5�X5���Fw8�J�''&�� .켷�(�Q�	�,����9Ws;.W���1��K�9&5E�,�ј��}��{�wY���&~+���G�H!͹��>ju��+n�a4_�̄w�����s&�&��'��u�x�~���-���@0�[����Ɗ�5P:bJ�LfJD���d�n���T���N\r6�?z5fԾ����רg����W�P�0�/Ϙ"�u����x��v�M��Z$H���lBxtw�J�r���K�M��1��<�1�U855�B5�Ue�Q'�7��{c�~@�6��@f_M��;��nM�&i�[)JW~�2(��z�oO�����rB������ܢ�mB<�hѷs�o�?D�!�����DϪ3��Y
{Ҝ���������	��_C��۵(�[��$0�?	^��R�T�uj��>�M�?Do֭�oÍW���%;�?B�wxdY�lo�|qT3���5��]<�R�~��sq��,
��o]]��5H�W�'=��3�3�ڄ4h��.����TtQsmaw�N�/[�s�+�L콣���� E��R&g���I�?�NI�_m��OK�:Ύ����D�+�$�lHY�<<�菮�e '^�NO1��/V�0O"����yၫ {��٤R�د����<�K���~�t�A�W-�i�i�-e�F�t��ϑa+�Y��X�	H8ƟW���݇�B��ZG +�Y�8� 8ߪE�{�xn]�[+�����c!����ƙj+Ʊ½v��0F2j��9��q�y�F���ɣ8F��#&�[�)l)��\F'`�j�-==}�+���yCaa!g�]�l�3�\~�����#V��W��EEE���.�m�x�R���&�U���;�/�p(%7�%���ӺaY��RGH��K��m��K�4�芨M����O#�uz1�c��;3Ir�n�R�L5��rnr6,zwZ�����ɧ�s���ׄ��F,���mhh�aMԝ�-���fo4˲��U�{K�+,���[�B�fgg3�j�Ǚ��m�/��	�\�<<b;v��N�g��'�+%��"q+:�ӹ���L�Է���s�g;!j�]�s�C��������58Ty��}�_�j�Фo.��w�k%w�41�iM�V�n����զe]Fg��������#=!��"�]ᠡ��X�Z��/�.ۮ���m$��c������(Z
5_�Z��wu�}��ZQ�C��{�N�����r2�����P��fF~p(AES�'Jς`^���i!ƃ��?�%$r���+�R�� $%�����h��5���Ԭ+���P�w��=���C��t.���ּ�&6N�vUD�c>J0wʂ�M�Wg6}j,�f�|6�u
�͞:���"Ӱ�<�-�Nɯ;��N�%P<P��.�B��Z�-��Ѭ D�o����	��y��6��4�D��a�iC	�Ncp۝����J��8Дc��6���eV0D��؃�y�s�?�{����V|�h3�-���t�v���$��Ӝ���6��ey�����%���^�v�q��V��S޼y�֢ڰ��3o�i 
�@M��|�-�P���t*�����)����a\(:����NBb�H�)��w"DQ���s��jP��rwK��������%>�r��L��z0�F��6�y�|�Gz#�%hf�0�Y�FJ9�y��Ǖ�����z�ޮ�%<z�8��4��)��:�����-�Se(�w��r�ՓO]�D%�,�����mp�p�U{#�EE��Y'�}����3X�x�C-?�4M�s���᎗q�X�?*ydEZ�f���_, $��������E�*;׳�7��7�y���~~_�F����Sc����T�N ��� ����Ӿ>`�X���'������J��TU����&�������k���(����}�&9{�.�'PK   6��X�v��3  �B     jsons/user_defined.json�[�n�F�A� 	F%Ծ�͖:3F����<FP��M�L:��N'����7ͥ/�"R�1��`�y�R�so�*�9\|�ã�r�_}�i�p4��y�g��1�+�eR�:����䭽)�=�6�t1x��"���-� )���/�$�S@pv���3 �?2��LO7������h����i�Y+#"�JD�(
�D�Z��<���+�������R�2��g{Q"(GZ*���1p1�ͮ��4;�b><�s�-o���vf?O�4}H��b0����y~������!����ߖ�Bv�/E
�У��<-=}���'�!c@%bD8��7����}�x|x�(��/3�����d�ר����&�M�o��]�F������C����6`m�� �c`���F�̀�`{L��E��؀�i#�l�W��E#�j���	��W+2�_��]Z ���KE~�E������ցZk]���J)��eyFE������?�wg�$���7\*�e:O�Y��V�ߖ+�+��m�f�e�n�,B��콸�f~Y>>��-�˳�6a�A�22Q�G��� g��i-��h�;y���V�	 ����:}]k�g�:�>���T�Ͽ?���tG�O��eU�׺��cPJG�WH1� L]D8�y�x�K�]��c��Qg5�98��Qt����H6m~�(��4�I$���+Ǒu�<��Y�x"����>�#�x�(��/��0��B�4�� ����_L�{H�*�)&����f}�*�\ࢻ�7g�
V�x���h��\�x��`Lw��?�y�2@��n�-VU��������>2�6�qwl�.;	�U�~��
v6x�ބ�h�q�&��Y���0���'��mvyR�]^���c\f�٥��!�H���eZ!�"�8J=�]
�1�
1��Ơ� i�)�f�Ӫ�f�s�E�2�8N@��HU����V�:�z���Z	��Xr�GB�5�l�V��R�1k
�]�SN���T��a:�R��'��}:���=T���sSz_fY�н2��O
=�����P����0q(�z'�_M�����2��|�B��4��O�S"�@IQ�8h❤���l���D6B<c(�4��F0o��R�r�gb�C{�0_�b��i��@&�у(��7܃�Qb��xh��܇V���B�P	����M���%����UU��	��r���1�|l�m��M�ɖ���_�y����kd�'En=p��|k!z��A"�(	�6H�H��$>c���|�;�:�sp�j)�R�Ȟ�AA4���)A��k��Y�F�pĭf� �9Ca2#��m�WG�/�'"tÅ�h!�����/�7=;��ߓv�+����s�~���������c�ՔnC
�n9����b�oO	�z2��6�����R��#Nzp��wك���,O��7p��F^����������ꘖ֧��r��0�Q!�޼]�$���������'��!>#���EЬ����p(�x�-O�eL�q���)�u M�И(ì��)�e�$W���Z^�4�]E�hj�������!L@*$�D�D�s�w+Mؤ�3[�����b�C�l��"�^֫|��r�& �||���IDhD���ztec���5���(����v@_��.>����C�\x0�X��ȗ�����|��tkS�٭uOEzB��]�
o��T̳�E��#� � �G�L�e��߆�6g�����LQ�0��fk����8���/|~����|>.�2���Oo�v8�ZW�E>�䨕ݔ�Dp�$�)���&H'�(�8�\֊�z��G�)�'0Ye�_�۲V�-)�G�Sq���=�+jƢ.u��Ɋ0�Gd_:��۟.^5W�j�Ny=�n������}�KE'XH�â�*�����v�I�N�-E���P�	�_u��/�V�)�z	ך@u�v=ƍ������]̖�l�V���?�͠UR�n���y�R�v�Ǽ����m��f�*���#�e}��pLj�;¶�+�p�t�=n@R��D�ᶑ�T�EX7�)i\Un����&h���ͤ�5AKv�m�Z�TGXӌZ�tGT݌Z��J����f�*�(�*�QkuiG�f��5q�uDmDZ�xGԖ�c5�KtDmf��]�#j3�XM�RQqӺ���I&�f9] ��(a:��=��b�X����Q�˩��ï�mj=x�ϳp��2|YyYyYyP������|0i~aW�wD>�D�	Æ9ĄP���"�<EZX,�\E�U1"$������q��Dq�(g��i ���@�r<_�]�p@���\P\)�Aj-Fj��4�]%f�]%vs5:6ZRZ�SC���K���v��J
���>�O��\��N/�ײ���d}e��vw)Y+`%A�@�a""l��^#b$1I4{�|z=�6Cl�-���}6�Hd��1�}D�CQbAN�����+f,IPG2���3*�M��fA��@"F�B�U�I8�-[O�ш=6B36"�ұ�Ͼ�<.�����+�"5��}�։�5мA�:���ϛ;�:+T�;����݁�	��߀W=
����ӓ�9~MU�o���Y�k
4���Z=�BK9�n��-�Ǻ��C~�:d�"�!�h.m��O����4�dj��� R�T@�*����|�	�*S����'�3�]B��B�0ҞSĩ>!����l�|��� ^j G����E��b�#�!�����-OQ��=&Q�^s�'��%�^s�\(u0h�� 3�(���3�B�兆��V_#��]/4hO��eP��5��SoC���=���PK   6��X��f�>  @�            ��    cirkitFile.jsonPK   6��XG�~��  � /           ���>  images/0739a1b1-a163-452a-a325-ab452d55b136.pngPK   6��X� ��! �3 /           ����  images/199a26a2-2ca8-4fec-b52d-fcf4e34cacf1.pngPK   6��X����7  �  /           ���! images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK   6��X��D>  ?>  /           ��&3 images/681693c6-5654-47c4-ac94-4786caa34b62.pngPK   6��X���&  �&  /           ���q images/6cd43c8a-9a35-40bc-b660-85b087cb5f0d.pngPK   6��Xd��  �   /           ���� images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK   6��X�1.:�  )  /           ���� images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.pngPK   6��X�Ƚ׌  �  /           ���� images/9185dcb2-65ea-4de0-8d42-42cedb1b5634.pngPK   6��X�&�}[  y`  /           ���� images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK   6��X?S��� 2� /           ��i< images/99226213-8268-43da-ade8-d9d07cfcec9f.pngPK   6��X	��#u } /           ��M images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK   6��X$�8�l  �  /           ���� images/aa130aff-16e6-4627-9689-819d55b5861f.pngPK   6��X���7z  �  /           ��v� images/be8de2bb-09ef-440a-a2d8-19619bf9d0dd.pngPK   6��X$7h�!  �!  /           ��=� images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK   6��X�GDU7� �� /           ���� images/d628d844-ce42-4e82-be63-f5fdfa438334.pngPK   6��X�G�#  �#  /           ��� images/e0d0e70e-96b7-4f7c-9039-c9e958c885ca.pngPK   6��X�N��C� ~� /           ���� images/e23486d3-0dae-4ef6-ae24-86700798fe45.pngPK   6��X��[*� �L /           ���� images/e5080447-3a09-4b80-90ec-33743b39ec87.pngPK   6��XP��/�  ǽ  /           ���d images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK   6��XF���?� Q� /           �� images/f590943e-678c-44eb-a174-3243ba5f3820.pngPK   6��X�v��3  �B             ���� jsons/user_defined.jsonPK      �  �   
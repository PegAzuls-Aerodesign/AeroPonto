PK   O�XH���
  AW     cirkitFile.json�[[o�8�+��e03�(Q~�vf���`t���D�֎"yd9i7�_RR۲M�5Z'ҹ���E'�SШS-��1��l��
L̃�j���?K�����m��ڨ�*X<�c�~_����2U�̴f�1CE$�"#id��L�$J"��^�`qs7�aq��8�⧄�0�y��X1	M�C�02�"U��e ,�8�N<�8q�O���"	Y��,�Hy$�{	>c�V`��I�i�2�`Ls�i�Ӏ2�0�)�4`LG(��d�2�ာ/�,0��0Ya��
3���;5�������0}.^��8��sm��̎0}>�'�C���:��)s�Ε���;´��ϻǧ�.�����v� ��Ax��;-��(Fh	��"�h��h��h�^�$~P�	�~�����q?j� ��A0�a�c؄�b5�A)W5���
��7�X�<��a�7	�FM���P*Qj���������db��O.�~r13O}�S&.������{j�9�L��=��x+O�/'������{m�7�j�-�̶mT�l��Z���EK�E��%�%��Ezђ�A�'��A/�_�����3?f~0�����A1�A1x��~P~P~P~P~P~P~P~P��������m1^�_���m1^˛�4�-�ky3�&��/Zl[\�om?+^�[����cј�r]�����F�&X�`�G�t�ws�_;Q�cZ��6�4�i�i�c9�ØF�YXpw�u���lةJ������-�q��h�{�J����{�Q��H�{�X���ۢ�͔v�u���Ӷ��q�9h��R޵a�胜2a�H�)#�%R>��	�G, �ݼ� B�E!�°�E%�,t�#}�R���a
g72:�bgGG����H�H��8`1X�6�6�6�rl������4�OMK�'EӢz��hZҙ<;¬����'������s�#u��^����V��5�S��^~tݡ��]�[}wCF�����ݟ�Y��8�ce��9f渙cg��9�$�I@��I�� 'N�8	p�$����k�S��m�����~]*ӺeY�oɎV��7m��� 9�� j�r&7���/�1�8���� 'w�̎ڒ���j�n\������*5���q���v�̍��#�1	�I| �1)H�$�����T��r�6F�V�T���,6m���Sv��E�ʞ{�N]7��4ma�zq�������m����R���Q���*�����5�j�Ua���ͪ~�T��z�E�ʍ�či��"-��\c������m��^Խ�����mc�K��yҏ�<x�^Y�7E�튾	etb W®�s��EL�"���BP�4#�BJd��X�a�`�[�/������VUY�hRy�uSX-��*h���֩/��4�ͼ�!���>h�@ݩ��I��i��\xA.� _�K��qz^��4qAgtAN^�K�˅l���1�Y�G��q|DO�@� Gt~DG��.�u}9�C�wk�r,���]ѓC��>]�.f��y^��4��.�o��m��ݴ��6�����) CM�	#0$5L�T&�ig���.k���ޗzY�ej��ĆkJB�"��̆��B暇����'�<�a�Ɩ�P�$�C �L��HR&wr����Β�I9���Qi�Z*�!�2��
s����P��8�ܾ��+y�*J��Yڴ�%

$�R�rIr�)8�Td@,�{�4u�im�=-��,1BmW�^Dq��4K�0:�P���ޘ}ot�rIgV��C�bDp&@��eT��뷵��qr.��s�����T�#�:��Ʌzh۪��{A�>�nڟ�n�f3О�lڼ��9��bP]���k����K�:��v%�.
M�2�^��� �7"+�AY�ٛa�ɉR2֑�S*�S �y�E�̉��PY�)Csb,^3�3�Lr`&�)�CJ�TX�%yL�1Q���S��`Yx<ԅ�mL�]��o����j6�駙57�^o��2sܳ�i�|�ֳf[�j[����{�t�ʺ>��^�	5�Y�]~�W�{�ٔ&k;�t^?��<��?]#w=*ӑ�Ѷ(�^��ۭ.�]����'Z�Ê� s�8�q����ǔfL��<I	�,'��ab�Y�ei���u�������_�|\�%�����Ԧ���8�J�G$C��$�t$����p�	�X�rs�qK'�g��;�8��΅��~�]��,�+��{�z�z[�mk۽D���^|�����S��nW���빕�z�E`��U���#�����Ee+�����ƴ��/�y��{K�=�<�б9����5����6�uQ��C�>�T���i3�NU�?�t���՟w뺨�kծ:]6m��y�S~������.n�w�]ϵ�C�=ts����
w\��+�g��y�u�4��{�����d��� ����3�"�(�C�� ��n�1����Y0N��{�1� ��N���@��X�@�+��� z-�� ��IhD?��?L��1�i ���|�{P�@�/� zm�ng|Pv�qu�� :�-����l�@ౄQ� �%�z �a�.Ar�8%?��'��י����@�c����f �@ϔg�,N�o:�@Ӹ�$ ��Ε0���'����<���@����Y㸥��%N�79(��S�Q��)Ti�6�A�_�?�j��w����ܻi�͝�ʺ��c���ɚb=L[���PK   ���X� ��! �3 /   images/199a26a2-2ca8-4fec-b52d-fcf4e34cacf1.pngd{eP\A��������݃���u��%�BBܝ �%�Kp�`����߭�����vg��������5�1���@ ����.��!��B�	���TwC/(���.��^�%�����7[o?O����������������	2��� ���a�A1��T=o!�Ŗٖ���A���GT噧cԅr�k��,����vH58Q�ͤq�������Å3x�HI^c�P�~Q{��gxei{�v�Jv�"�����pI��í�m��͔	��8�g� ��v)�Ep+uc�aʪ�b	D���� O��8x��A������#�֟���OQ<#�����F�[�<Q�kU_,j	����},��php��E�l�z���:^)�����z�o�FR"��:���y���B�	��.���'�җ9����l�휗9d	>��z�w�/s��#�Ү?��@��C�]��s9�����D�z>�RF!�Xj��h�G��rѩg[xq�h��2�i�����$id&�`EQ��R,楚�Pĩ�W^ }��ƽ܅c��??���`.q���d���/*�
�9S���L�(���{���8��j��ѹ���b��Mҥ�����U��#I���ջlA���G�,��ϐH)l��̑�������Ļ����Ĳ!��jV�H��`bG�ϻ�2.q�",̮����H���r��1#��OVp5�-A�[��%��q���H��]���<9�6��&EB�(R���n"0��_�մ�9Z	b�@���&�ghk����������.n��x�}Z�V����!���UT8���<<
]�`����s�ǔ���{��x:_�7�K�!���B��Q:9ځ�)��+Gг����蒖t��d�E+�^4j-���?�|b઺=hzQ�w��)!�nա�9��
�-�W�_kVg��Qe��7et�R����edע�g���T��{T�q�O/dՐ>�o����5c�,�����}xW�$x�)o��_���ƈ�8�2�z�#��7~hP��4�h��}�/���'z������و��ޟ^r���}pCY�E��~� �p�J���Q��[�y�f��� q�+FO)#�$���9)�Y�����������o�*�*�����]�{�3���Ji�<�e�y:ɣ{��U4�bf��߮	͛ͮ��e�i�<�#����~g��Ro(�8�EA�{�`��A�������ټ6JńY�-+��+��ȤX��o֚˙���6�J��}�	�`B>B:�_uI*	�����VB_@�q��������r�����l�����7�t�<�D�ë�uD�Hw��jjǢCS����t�H[`}KL�O�38����݇���R@AzE�h�"��n�T��Iy�.���.���^y
?ܲ��f�;�i�3SU�N�Ä��	��{J��� �z�@�������[s}{]�,�i+E`ЙV�:�y����ïH��wy{)N�o;���^<l�~Ic�
�������w�Z=%�^�X	�ů���NWD
�j�d<�N-ۮl�
{E��������|����=���?}�"�$� ��#���(�vG"����
��P��?D�zr ��j���`�����l��0e�z}�~X��q��S�i�Qʸ���A��a%�;>�l�5EG`���ul$��̍#�EOC5�G�>}�Br�0��8�"=L�o�]x'�^���wxz��~�S���.��NA�d���Z�p�~4��Y-Ƕ��=�L��q�̸WO�s�*{���Qf�)%��H�¤��:���� �K25��eË�%y��@q���	K�"�ŗ�c�/���4���oxY�[�	ت���"}?>�eF2��(*8�@&	|���%/��b��$�m�
@V"�83�`Q�������c��D��Fx^,g�WeN�R^M6Ŷl �j&O�DE�^���� ʍ�G����s��Ʋq��r��xVa�*x=�^�pEt}��҂���k�$/�� �K+��v?I��$iߞU�M���2�;�;q�1��b$��a�,��[څ�f[c�Q��Ř�(�c�����ڲw!&/c�3�������Tm�㉗����nW��7����-��r瓚'!�`B���
���>Pb�a!�������M���p���u/pz��Ӵ�s�'L&2�&�R�MY?� ���B�֞>/̂+�]�����`�R<va�LZȟi�*i=���)z����ē1|Y�D�"�QA =�3�`�2�b-�����r�/Y-	G��tk+h����^&Z�b3�I��/�M�@}uf/�ሺ��:�b�Y��x����ǳ��զۭ�^`��<II�L<�ۖ@��z>wD�:I$1((��{������}7�.6鯿��XdYX��J�;���h����0�1LO�78
�����������5u	T-���?�œ���Z����Ya:r%��<��W�S���i��e�0�s9�hi��I�)���OU��t�u���6x���zA���}��l����d	�1��ˀ��7��^����S?�ʺk��O�bG�����3{����⬰�pQ��Z��'�7�s����J���=������m����$�Nrca��Bn����٦4�cЅ�(�nTTACz�� bg�ϠU)�n�2�g�kƹ$��_�ߠM͞��T�u��R}>!�s�U:��9�����y�QQtLEc�wT+,����W��s�7��4v%:#JmiD�ٕr�2��S˲$�U���E����5�C�e+2���B�&��P�?8q�ʘk�`�0m&9����9Ë�Zﬀe'P{Џ>�N~y�aܑ�,���h�>��cY��E-�D�x�'�Нv�O	�T�u-Q ��$�(Q�4-ZI��ړKI�J�ײ��Jr���.j�Z�L�#~%�J�s��&fEyq��yjB��?rO}�i2��������Fz��_o��(ŠId2;�P����q��@�Z2&�ؓj�F�^	s-��u���^ �xG.?��d�5���W��+�|��-�^�%{92'��z���K]V��O{ou1�N� *�,
�0~Ca�(%�?��-fx��*�b�= ��i�<M��Kc�z�J��b�'���Mw�d�3�*@�&G�_��*jW\�:�W�z�"��hF&�--�^�6:p�S������ͫ�N։��KL����L���e�R���2�� �GǸKǵ�^�^ u�H���EJ�#�����V*�	�g�m�����9���"\-���%��d�/���#�F#ˋ[6����t秫�wf�ӮTF�ߟ���+�G����H�`�mW�9�X+:�K�25풮���_���8�a�
&�G0�Ac��.hP5�_X�Y���b��]��0�޳	�K�#a�54K'�
 ǂj-F�}�z�
�totIo�/y����b��5��!�h��T��D�������N�݌�r����ԛYOʸRnIJ�ym�-���g�:�n�I��.WU6E���;m������6����T=Wb1igG�ԍ�~�h�8���}�����D+	�#���Z3	�w͒��U�^Hc ?�jn��p ��|#������% d7$�Ю*ǝ��4\)V?TP��PbW�mN<���'ؑH�ZbջH��,�i�����!�����]���� �c�3*��Z���tG���pؐ33dS��Tу���1��s~�>fd���+�	����_�ӓc��?�.���b��УA��;+�����I���J<��am'La�l��������;���dͶ�!u���
x�]��=sSq�UVi�Qb_�M3��Fv��t�6�J�Fv-���fki�B�('�Y�FJà��s�kiW���P[�p?4		�Y9��.������֙x>>V1�0`���TNLSd��y�0����!��#�v0��E��%<TK��,C��z$�6�}�����V��A
W���y��P���������W�G�2'r������Я!�Xǎb���o�Wﻈ��1FZWi�\�Q��_Κ��JFQ�{�׻�:Q�܋�>�?ny�"*�U��#��?��r�FJ7Q�D6z��5���()��E*��708�J�}?	�`:�O�4�4}��1�� �F����]�@�Lͣ�L��ۊh�����|��F�4��ݥ�����O-����-��誰��!��vOr;͇���1�0�o� -:�l��\d!���+'֗O)���wͰ$�L�S��Z�,��/`���@��{�@@bA���9]��q� ����Bˁ�7UeݭQ�YG���s��=�J������GN�w.�E%/���v��/����hʡ[�"Ek՞����Nt�`�
D�������H!�GO����S�	;�UP��t8b� cL�A�=MG���' ��T��-KH��KG���:)e3Y����������Xw��mĆ�����x~�����<���l����M�}��\�`�i+��M�gzu�]�ՀA<��Ԣ���O��4L��⏢����cɋ��7�$_%���W�
��n~Jh�/:H����|�')7?���'@�|JR侄)L;����R隭�����0�/��n���W�E�ܢ��&�E���{�Oo��|d��MM��'����\���c�H�#�c���?<�2�Ua(���}^��"����>֫�����U�k�nK��l&�K�ۏ�F�2�fc��$Ǿi@}�c܇��.��)��I᥃��И�a�s�-������ƿ0���9��ó��_7e �rſ���!����U� Ds0E��X)e��i���-�8�b��O�؅~�1"Be%ݼlD�\^��|�4��E#���є��uV��"f�_da>���3�!�8������|D��_;l�"Ҟ|�>{z��m����I���i#�(Mx=�5��рA�Dq��?����7�y~.��C�����!�j�q=]O~��^�}��-�L��eaI ��.����{��sH}aB~"�r(t��=fW��u}�z�{f����t�΀F��r�ZHWtB>s�i��#�b~�L,z3ܶ�|31Y'�x�k�:m͕Niɩ��)�f������O�3��o���I�"T[�J$���~U�oh�B\�Vx���X�����LK�����T���'���V�o]���܂�ECM0-zS�d��EM��c��â��n�U�A���]�J�w�sg�C�}��P$l��:�n������U^Z��P���&���o�-��w�6���W�Y�Z����|�jU<W�|r��:,�B8!vcբ�v�#�		�d�a���)pۢ��񟔡�_1B�&~���e�shF��.�®+��!|B�y������R����/4�L~Ws�fЅY=��3x�/��t������߇@_��kv���{�����@X�˟|���H��1����
w��#��ݼ1f���Đ�dv|i��47%x�������A���a�=�K�E��\���Y�?�m»��A��ju��Y�eD�vE�~���&�1�ްXڏ{�s�tD�y�ῗu�mK-z��廪��ɛ���L���2�fd���Zb=3^J�!����Lzc����#���	C@�B:��η�Z#q6�T\Z����M�f�Z��υ��nd#YX�$�󀾣��V1Moa�<PB.o��^����%T^�ڣ�JVSmC��P4�*��󒿌�^9A��Jbw^�6�滚����]��M������4��A��S�y�)��.�����j�+֌�2M��*L���X��_K�|&;�^V<��,�~cͻ^�}�߇����53��P�ճ�Ɩ�E;�8����Sr�KJX�\����.-g����i�4��Tp�"��@�M��)K��mR��(���I�>��]ރ7��?z�>8T��a�N}~���HU�Jh�WX�a��LV�C�-Q+&w���x\����[��b���=|nu[IFӒ�����g�q|/�n��G�^�	X<|�b��o�w��n�'��8llC�h�����I�� #�Q���`�����Ev�y�̫�=��v~uRBu�-\z�$�zf'!�ی�KP?rZ�J�앯�w���k����yH��'��K��Eќ�G�H����@'��#&�����'�R�.��Lb��(1���)79�aq�!d���`!�m��<��S�ו5�dO-�E��\��P��4:��O~e��^�͏�Z����x�pW�]��p���B	������-�%V�*�z���w�����iiy��{�Q�'�c'*���W`2F~�w�]s��`��? ��8��+���#����~GԷ�L����fm�ݝ�e���C�[��4�_�����0/�Fxu�<j�������Tw�Rf^��i`4f$ ʎ)��px�CNW�)�'����"6� Y�� �P~�,�,����Ik|���I�0]�5 ��҈��t�d�d��m���<�q���C9�k&���;v��K
�Di��	o��Ĕ�;"t�̥��߆��`D6�GB�R��g#?���0-���%M���c����8N�+I���FH�8��M���QGr��1�9���M&4�|��<1\Ƴ��S?};�(T�QRմ��������Kj�<UT��w.9��Ƃ��W]|s���մ�`�ѣ�ܨ��IB�}o9��}+wa ���)A&e"��S�f]^}ɸ�'�i����kw��4��Sek�L\�_1W6t�Bo��_E�X���~'����=���>d��$�C����т��uj?�KOԬw��Q=�I�H�)����4��k�Snc?����0W:)D�Us����.���T���L�Ј��א_�`�x�9U��*��?ކ�n'xe.�H��IbG�bV�Y��bw%2�`ǝ1�F�ڷ�����QKV�
{xd���ț���Z�<���\5�����oY�\RWry���J�UT �5���X�EE�	�ӫ ��C��d�� v�?�k�%T�bu�����ܪ�� ��*E�4��ߑ�]�dIPۥ_N��X�񸓼�n8��6��7�K�j[�G�B�]T�W��N:�}�[�*�1�;����Y3�;��.�Ru뀟�"��~-3:�ug<��g�L�#�I������r�C��"�<�z'��뙼�ET�(g�hP;\�8�q�͵��9 �%!�Y�O�����W�I�0+�"C�v���]�K[KLܽY�h	ie� ejf�He��������[�C��]E�� �99�>#ۍ\���tq��fW�#�������p;�[?蟓XmA;F����awjM��w�A���+t��!���Y���nץnt�!�1�b7U��c��.��<պy6�)��3�giQ
���T���+��k���J�v� ��[���Iǌ���!�N{���zQV��%L��^������@�t����|1��� ~a�}u�)��1nt=��2�#��N���6�9������Q�IDK��\��������Pǭt�η��}��v$�_�[^v�bFKk�Ƹ($���ͧ��e�'�6�x_��9�F�ږ���,/IBI;�lQB�N>@�U�ȟn�i	il�mOL���#u.��[�^����:��$!���^�q�䭭Er@U�P�+fʡ�/��Ao5Y���	2�����p�Y8
c�#ؼ}�h֙�bH&�p��ޢ-���O-Ufs�G���-{�8�M���c}"T�d���} 6V���M��u��H���Y�=13~�����*�Qyu�v.���Կˋ���T����D�����C�ώ��ꂴR���>���c��]7/�e��9��L�g�
Z��1�h$�q���V}1�60f���I�ۃ�=37}����E�vtT�W��Lj[�HY6��f�cG��f��=x$H�La��ub����.���y�FLR�|�N-=��v��_T~?q'��9GnJT�޲}��D$��m�rb������v3149�(w��ܩiyV������Y��P���)��RĮ��*V��[��_7i���8E揷�ڦ��$���(�@{l�"Z�]�#_'9�lO�o�cж�T������gs�)�LH<ұ�����g�����"X�,��Z���E������|��ղK��0�}	�17^�z���mVq�!��?]��W��2�rhT��Ր#�`W6��TX�Ҧ��mZ��ƅ���cn��Վ�<��O���r�|-��,[�,
6Hˠ
�#�|HN�w��W����(>�-H��{��c�%L~(�+��J+��r��96+(�	���hל6ͪp�H�{��{�8��E��B\_(����t�*{n�6�ݫ���
91˵7�Z���E�6����ܦ�?g��՞��j���PY]�~��_@��囬���̒�<M�{D5��{����J���[� �!��7��񛔏�c�ba��}N�)�����j�G鶬�1S�٬L�a�%Ҙ�Ť����\)@����4��������lV؍��m� �E�"9/�K��b�eC��K�qw�t��}$�W����g��{�����;����x_��'kf}�u��e����1�U�篆�k�7�|<�+j</�I)����P>d\�����	����ڧ4Eq�xvW���l�t(�z�:�H��=j����Nf̉��F�F��͇��o�!C��q�" �'�����4�5�[S����w+)�=o�ܔZ;
�9�Y�Q���G3����W��a�PV�	�@%�z- ����&¾�gb���*g�i�'���$#�i����_�J�|�u�;��r;�T��G�q�u!p[���v0���ܴo�%5�8P�L! f�k��z)|���o4c��c?YP
^����M�EHg7�o�07y_���2Ƕ��Lj�w�S��m�0�_�Xk��DǴ+��v�
���m�KO�<S����U�_�o�3i�FP2eO"\絴Ay���0���4�86y��QW3	���J�s�zY�����8*TX�������0=MG����(��(#R�q����a,���(��۞�}�0��6�wC�ߖ��0�F[���(��ٹ����b�'���j�[�y��k>���Q5��mqVE)��:!sC�[�3ʸ�_�4u��K������(�C���`j�V�
�����J�4�������<~�O뾋�cl�v�Xt�N���~Rn?���`�
�RjHV%Mu�+"�2�����d�K�r�eF�)A����nL�5d6��q���m��ʿ`:����N�g@Q�nqF��J��}2,�-p���F�.�t����^�@B�����A3(�������j�6���@��v��#�Ƚ1�T��P�J�q�a�	Rh@�k!��mNR��*�V���Ns#�;5T�K��Fd����b`>]٨(��5��T�*����;���Դ��.�V������:����#����vO�1C�M͗���1�%R_�O"q��;(G�J�5���c�y�1
"�ԑ�K3���]"�F��1��gM�f����E����[^[������xݾ�z]4�n��������enNB�>'!���KԢ3��n�5v��#~�L��aJ��������R���5�[�^��Ư#yJ%փ��[���=[9
��;�i&���赏(��>p��,�]vV(����DV�kC_w]&�!��.p�8��8`��-Q��vũA<⢨Ǻ����o�m����=�?�~f��2o�+Ĳ5�ب>��`*K��~��X���m;�ʷ��n��Ն�6w̩���a���&e(�~��s���KWf��0��ϧ�RK&�2�i!�zڊ�ay�H���\�R5k�Tc���Ц^	",�,�h<�0�7�����}�~/���Z��H&)��5�IY�
��� �hDY�F�E� ��;�m��`1��⌳%�i���o4}x~�Ti�2.�)D/�]�U"��(8 -�}�\5v���i������:�80�,Z����	�+oXJ�Rs'$�;$?BE�i��y\�ZL���ۿ�������sn%9>�^����p���kt�����M��'�₳���T:�~R�Jz`'$ŏ/����S�	�9���=�{*a��+Sd2���S�Bbmc�q�	�/���*����k�x5��%_V�>Ӱ/-�n��#�ɠ�R�W�6�����23�9�l���N�e}x���E�˱\�,��K]����YG!Ʀ��آ
S�xu�H�-Ȫ*�!7�L�����^��
��xS���PEl�Di�
�L$v�N@���592���$%EKEIדi nxC�pϯG�~U0�)�"�me뫪���T�2=F^|������Pl�������)$�^�!68XL���!]���N}\�j����"���0qb��T��K";�?�����E��Q�l��DĲ'�pމ���v�*zH�n�R8k���n.e����%3O�(��]�K$�8���`���@��X�嘯���=v(�44��3�<�q6��?���]�:�M�����#�(�_q��0"�p\����+Q׷h)�"�
Jf�Dr�B���J�Q����x]2U�zUO5��s�
���v�̣6��m��5%>�BA�m�ه0�*�pe��e4-Ҥ���RW�U?�DN�F*:U$󎜠��(�?aj/rG��dۊ���)�Ψ,w'D��;��Kga�i_/K'Vx�A̪R�����9��J8���Cj�]�^����|q|�����N��5�}�&@/�M�"M�>Y���]�Z�
�V�ZU�A��u䔖w$�$sS虳'�/C@�s-�ȣ0p�Ԋ�H�6�q��ǩI 6���QW���"�	r;�}�9�ϰ����(V[�YG�RZ�K|���%~?Ib����@�*M���㊭�3�iz�]"��:V�q\J�����al�t:|>�8��V��A�u��<�$�q����@ۺ�
��9����ީڈ֐��OQ�~&����?!Kۛ�0zg�)�n����`�Oa��
��n�O��}��B�?6c��G�8���1�}@������!�9E�e����|�4
$ݲY��j�D��I��@��K:ڱ��0�5?F�}|�����#�k�a �p��x�;d�z�<Qf�O;J�| Qj�
n�=�kOj��.���[8Yr���(��3��&L��Я�_�_t���T��L>�rR��'���ӫ�몢�4`>Ja/�GuI�A����B�S��!
��!2wK��%�,!q�ag�)e.������׆@�}չ�T�nY�a����7��oUVGl�ӱr>^�T:���O��8=/� �78�{׏P���:�^i�K��u�`޼�*[�*�����t6x��d��\�WQ��0��x4TB�C�P��[*�Ph0�_���o�g�@4NE��*�:!��6�=pVLp;�����i#9�!RB���!�a�lx�g��Hf���J¹�8����L�e�ƨ���i�D�$��gQ��r� b/\�8b�-��)�.�!Yޑb�~�Do����3��?�Qhّ� �' �a�t$l-���-��HB�R��T��*'�p,�^�]��Θt:��-B�rroMd���s�rãx'�~F���`�S�"��͠���)#L�?%�!��E�E��Y@�)�<��m�-:���>E�z���̩�N#���A�ސ\X�-�KBTga#$���V�����f3���Sd64}�v�k
�29�QSҢi��e�:z��B惛���ՔOi��

Csl��9XI\-��̧N���e��1�-�oZ����A�Td���7�+��0zYn�/c���&�48g%M�X����jԄ���=ƱR��d���ypS��zHd���+r��Ƒ�̏��|fƍ}�du�~}c���&q�sZO���G���7
���S#t'�:�ہ<ǡ���-�f����8�!�	x�\H�<��0U$Y[���8�k&��z����գnY��R��n�f�Kjv��wh����b���֏����(��/0[PB�)���%>��i|j��BJ�k�sM͹���v����Nj�s�/��68�b��*ѱ�!L���Bt�}iZ��n���J�W����v�|��㏁���K�"E�M�LT�5**��������]����;<yVC�!�����7�;�@&'�v��s �U�7���9�EI'Vj
+!HUYZ_�$���/��:��`���[�~�MU��U��K���f�e��vO�!S��/�N��6܋s2���X�z�:���͚��3e�':�2)��My�y�<31�� x�N��g>�5�5�v&��_c���0n����4���4?i��L�L@��\���	`O+̙��H����B� !��m2ݱ߈Ǧx]��X�Ô��QA8Xd�d��g��w#���޾(Z�IP'��ܕ�Y��՞cv
�A�yq\���
� �wb��=�L�I��y� ֩��e�� ����
A�3r���"��S��j���
�����W�9%B���^Y�鵏�Sq�HHO�����Zx�Z��C��I���D �͈E_l�S=�=Sx�>cp��|�h�®�D[�=9!K8]Y�F�� I�-M����\u��8�h�wЯ��B�|���ɭ���D�ˉ@ 
�3f�����1(mO@�ĥ�����ئ��@q0����E`1���T���L��qK��`\��/}���^n�` ���i��8BO�9��Ht���m��%^�^ݍ���j,"�	�+�C1�� ��~4���J����D��Rrʋ�{XM8(�f��|W��X<�ߎ�N�J>��R^"d�rn�n��;3��(ʞ�Cy�K2�Z7�I ���#�c�L�g`��#�kݽ}�`o����#�G\)Ξ���"�������'� �j�G���S�_P�#����.q<Z���џ�Z���dȰ9�	��n.�k��w�%�sYn�~�-Xrs��j�M����e��A&�Q��1f�M?�=�J�� p)��9���IV(�b�J/?�mŮ�J�6�iҒY�g^��	�/:z�;{g�74���æ�q��ӼtY��4��hϭaI�1��řD;w����?��a,۷�V�,�ݞ:�;�q4�T/}�X���Q�+`?�QgdoJ ����_�Y��>/স�Ce��iդ�����0��n΍i���ز��m�*�UQ����q('[����|Ӄ�f��L>��]�J,��3I���S��fN4�Q�<M�A��[���V�����L^|��� M~-˩b�6�`�ɾk��R
9VE����a�9�,s:���H29ֶvP���0>���ۮ+�s���;�ͳ��]�Ԋx6�<_Ƥf�
���-��eu֊%������?�A\j۷_��K���D2��W��.�5a��%EII�]���	�u��l����xO�{�|�KM���ۤ��A�>V����h؄Գ��Q�r��uq���`�n����]�g���_G����������<5��ޑ3	�(��o��G���(�uS9� �����v���iY.f�C�Z��z��h�=��4�/!|$Y|�\1�l_�+!��I�lp���]j� U,���E<z��y�P���}c_��Xo��"��R��"Ķ~���,}�J�ː�k�nl��f	7����-E6mN)P������$ F�(L*v�T���w���0g�[/��U�E��h\�y؟R�Ս*w�T��������};+zF��<���JBMޛ|S;5���f򥟈CFnCH�)8؋	\��&X8k� Bk���l�ec5�{�r���{Qek�hf��-!҃t %1,9/�ڈ�{}�6T�!I���JxY�C�����>�����ֱ�sts�遌
�H�c�5���I6�c���G*t�lRՀ����q1�d��*�:���ⱈwG�2�ȯ��D&��Bs��Ӷ� @��E�����\�?�F��w���qNN�R��>��F5ل��<�|8�Ve�fHK�1�:Ǵ�X��"j��y�����B�k��&���_�(�xAE�,��NC�䞫02��|w3�;�Zg"�Ժ��kQ� 8���xA���J��=�O���Ob�zst�2���4<�ӧ�v�VH��3E듫¸���&����=���[S���f��an�-��We"|0�6S��'k��oJ!}E�I�$3w/�Ŵ���t�a�;U�?��Y/c"���4�N��op[��~^�s[�����n�8D�)�mNߍ)�9:X��Y�Q0kC9[MT��f�*���;�joUTQ����W�X���8p��'0�$˫%�d	R_��<��6��c��\)�l�I3gn�(tf��!
��j�jI��(�~��4���]����S�)�"WZak�a�|�����Uv���'������c�(�CKNP�/�[�;��ə�5�@i�Y��'�F�{]�7Y���l��������\I����!�N�L(��̥l!ϫZ�W���;�@K#L����7]k\�2Q��$�y��sZ �ȅ��Ϲೃ�Kk������ҊSk���c*qa�U�j9n��ϖ��=P�u��b~5�[�@+X��|�|ۡm� qx�r�e;�<��������o	�+�:1Ӽ�ӝ��MS`]ڹ|�u��FB��+��)���7�C)�����q�K͵17?��X�I����[����䭣���]L��k+��M�'Hf��"���Yq���Y��/�6q.�����E�*;K�LJ���߸�x�o��u[8���<X�*{��H��J�.����=wq�7Ҫm���h�Q�(`���k�@n��i{5�n\����[�Kfa7lg� �MVU�L�ʺP#ޫ~xz����e:�����)��w�f�Xd�{�֍C�߆6��i9�-I�te�fl��� ���0��G1����A�L��H~�0�V7��޽a��G�s�Z?��Js�	�i:0�&\�{�~s�i���d'���ī�m���?�2�8���K����O,B����q�)K�|�Dv����Vsd�w�"���]�u�26u$iO�,�y*p����n�݈�b/���p�ݛ��µҎ5�Q�d��V4��D���b;�9�E��痤נM|]9@:V�E>��S,>�x�	��&]���C��8�dǑ���|P��`+?@�1��S�Ԑ���`۳�6��/�����wQ�5B�p�-T�q�;â��d����yս؂Ui$�)V(1A}4=����.�,{���t�ƭ����%�Н��g	~�L��	��+�^�9�ןo.p1��@C�*�b$��ς��B;�ՙt��7�G�G�ϭb���/����3����z���@�&��\���"��"/`*Q��Dy�]�艐�·�M-u.c1���ԁY���v��P��0��	�ID�j��SD���	��zy����
JY�!�v�#$��֝;�5�Gb�~V�{�����,�{w�s�].��>M}�e|]I�h�\���i��9{ ����-���!S�g����'}Er@�^��*6௯)� �vO�/��S��S����d,s�bt �&yc�hH&$�h�,��t�=���R�y{���f%�m�fh����=k�z�wH�W�F�@�w�,����/J]0�۩��GP���*,R�Ϗ�G��I�����9�`,��Ѓ��E��Ϥĳy�gn�؏���+³{��T��޹#b?�� K1Ж��.!����|7Ϙ598�[r9�yU�꺁�џ�54�L���݇u�I۱�<	n�6DR$5X=.�>��� �4�Au��懎|��V�+.�s��6t�D��,�p�@��C2�bj�C@��(����`����y Y1���eim_g&&0��w*V鞐�?���_Y��QsZ6��|�T��u��_3�_�K]x�G$�g6�8g��몎ݯ�#�J|�.̯�Ԕ�&������X��cn�'[�G��J�N���J[6���_�$Lo�>1�J�;���[�/�$��ZL5��
�O�,��RP�+�s��y���y���9z�lVr�G)O�T;�B��%BOM"O�n���N6V㈮��d��&�k[b`d�����ǳ�v��B��Y[��5՟Ȑ�ˉR�2�E��U}d��	�8@	i����2��B�N[I���=a���$���S���.�W_������b��jֈsb�]_]����f�s�Ur�dr=����³S�k`D�\~B���Y	����Hǜ	ъ���aL�s���#-褕�k��%H�Խ&%��I���#�K�
U;t��Ŝu��*5�<N��r+D$C=�������y���z?�#dP)Μq�K���J�8��n��ə�N�4�������5�5Ì䉏 8ž���n�o���ܕ�	6R���� ����~|	��C)š:~�����5��Uۭ&QqZ}���8#k�;0�H��������C*�ﲾ�CfQ�vkC����"�gY�����[�E���CI�� "  �4�"��"��(% !�]R���H�8�H=�5���;�}�s}����y��b��^�Y�z���g��'���0��f���:w�tg$�	fV��?8�q^p�/^�f�ym�!����/K�h����-�*���^]�l�q>�Rܲ�����a�I�¡|dKT����������)GQ�'Z�X�
�aY5��Y���QV(}˝�{�5)#�	���k����E������O΅ì,V��F���	[^<�[=͒a��ǜ�x}�O>��̞���}�y+���_i���� xI�8�Of^�=��R�#����ƛ��G�9dD�7`��z�4��8�3P�!�Nxވ��/R�>S����+$�� �.ġo?<�W%	ݘ؝�~|�q~*f������p�Ʊ�Js�M�s�4��W��\�+7B��xc��婙���3J1�����=ϩ<��͍��,�!
M)�'-���}���zu�9�?*�q�x_��D�.�R�A.-7�$��F�]�CU�� ��j�&B�C�ӓ@0J7P�=�+y�M�����I�گ��>5������sx���������;տ\-�"@�k]&�^���!W��Aa]��F*�]O��T�����:�����ٓ�����k��4�}�
�r�r�zT�G��/�d�����WO�i���~��|�<�v�l�?�-����w+�i�]�=^�Y�Ԕ؂`��_��_�<�<���Kq�����>�dm���h�C!�u��/6���gM�Y������`��������}�*G�.�|��~&��u?�MG�R�����J��#x�z��+kF���k(E��<o���_�:��x�智�e��ҋ�����������i�N��g��.�p4|����g�C8y��m��k\��oK���wAB�<�Ql���׻h�3
�����f�3I\�����DLǌc&���:�>7i����	�O>�i��9q�A��Z��m�j��ǴRѶ�$M�>��7�'\�V�4sW�-��!.Fx�.B3g/���~��d��[��!���9�cZE��:RC��8�o?~ӽ�����s��g8��C�[�2�4V'����u�i��.�\)��L7;±!3J�>�jU&��^��=$i��Lw5�_��;����qr��s#u��]�m���"��U����^�_�mb.P����������+Gh�;�%�L���Iy�^Ȉ�v�<�Bh����~����諴\�y���܇��a(*nrc"i+���2N����mځ�	��;���q��^�i5G	ߖ����i�A0����1�������;�>�^^<���G��x�
6kZn6����E�}^����H�P�>r�@f�
;D�gԕ�9�>�dL��#Q�xN���h���W�%e2[�'�>,�g,��
J;�ӘG��?}r�N��0�AR@�Pa"����)�)���/�*ve�P���2w]�>ؙ���]4�M�}y��?�e�W��{���$�9^�8+P58Ny�>��8�j�t������s��JR��I[�����E�w�^��DA�`�v��p��Nwb2��P�����?I��=�ťxwf�}����eTA^�T�7������q���33����x�Y2�� +��-V�aՇ$_p~*5�e���uw4p~~�_v� 3d��B�pPk�%�\��T�<����yL�0�J���]�L,��zDH�ʚN�`�'�G�Jc���IF��3���x2�+�l�`#�~P����U�E�'_OeT��O��A��ʬ@1����A~�'�I�f
!�n!Wt:w�c�|7��3�!�+
�z(sRH��sS�>~Od����x��d�����su����\�/��f,)�ψŉ�H�*��o�u2l����������Ē����u�x�9xe^_Z�W<#�S>�{�G�7`�_f3��ə1�+_��b�]�7������~��L����`�9��[x��Fő`���ٸ�I"W�p!�gx�Q��=�Bd�~�퍻����|�t�,��G��fV:+��*}�U�=?�!�<�	l՛����BaQ���H�Wrи�bd�<e��ٰ�>d�Pr�q���}JdΣ�w���D��C�q������z�~������.?�x�<U��[�W3|6W�RCX>+8�I�ֳ���b��Bw�^�$�Ѯ�t���7yQ����������*��1�5x72
����v��w��;SN3����}R�*]�Е�ӳ���+z2g����E������׫(�`�kg���+�"���0u��%ٺ�u[Qˡ��ʳ0*���j���_�A��'�|_�~�1x�Z����R���U��|`��>u�Z8J2�񙸛U�/��^��ޝw�<kmN{�!����òؑ�<X/.�����,'+�B�P6�佺ƈ�������sm�@~5LL�ި���/>�5�	����a�Z�Ltlg����"����k�5*�R!�����*oK)a��(��ߨ8��F�����7{;ڽ��s��I��m�֚�XݹO�uwv���~N(hμ>k��+5d�[�͋��,˫�����!Z�f�RK�����H��J�ӣqVvȗ|��ɦ���Y
���1��yʭ����hH_�>V[�<P7���a1��a�����.wIN�����'e�T�N1"�<�&�Gz�Zc�=��6��Rm�N~��,-}t�M�ҙSt|].�5������=�I�7�!��:;;nWD6b��n��gh�c��3����3�W��lCms{!r7�Y)Ũ��mZ��n�d:�������a���Y��>��풹�ϪvQ~zaG��^�!qe�[���O�uy?�2�� �?�8tx�E�+��xK� ;)q޻��GhgX�ͫ���0��~��f>�WT���s��	z/,���[�߳}�v]���X�̟�0p�ZW񁏦Mχ�Q��}�n�B���|��K�f@|��L^.�zά��Ҭs���*������yO����02��%�$R&F���
}*���F�q��2���lr/.T�;y ���:�Q͗�϶|��R��xRn?749_��+;�Rϒ��A=��1w���.����)4،���8��fC��r.�uи��$JX-"��oKY�mn���{�=��A�qͅn��"ԙ��l��*i��:��D�4������Q�5ߍi������n���h[�@��O��Δ}wĖm�`_m��f����V`h�������C�����w8�n|̽J���.6-����y?L�8�m�?3e�9g�H>u��|�H���R�~�{���4��18p��dC����V(,��-32�xZ���p����o�2���IB�I���庂�+�:�4�OPO�
�Ŕ&�>pV���*�L�FyZ-g�Vg���F4�"uTD��觳���ԥ^i��M1��<�d�,u$o�g����Gh�_ ��7ܭ���Y��8�0Ezܾ8o��)���b�W��}�k�j{�L����H��ݨ�{�Q�kˇąuII���
���[���Wδ�5B���G)V
���O�fs� �2��[���m�@<����u�DK.Y�����&j�s��=��d(.�/�yA��.��V�X�Ϙ����+j��]vv~UȜϫ�0�D�{����p�������
*�=,F
�'p�X�I7�9�A��^�R�P��y�f��vך��Tp�u:�Ή'=]s	�T�Uߢך~]1�F��5�Ԛ�tC��l��/�߄�+FL��~Մ&�3�3�IM�y�*��V<�[J�$Pa�Í2MW��j�����Q®=��R�	��1��_Y&";T*ag���Ψ�4����㠒�eq��?E�V
憝&�%�x���Jx�,��"gv>��-�=>��[M�zHw(�V�\8��q�ҽp� �i2�����.U��<i�%7� �y����=GM��3�.��MA6�F���H1u�b�z��W��a��r�FT��9s�w��z�X9�A��������j`f��M�؈��
SuY���l��!�܆V��wLl�2ڙ�c6ɓ�9�̹�6@��*�L���Βk�z�=��:���n\��a�<٭:*]�<�G�[0�*����S�R'�:�^�����2��㊾�����l5�/��N�y�X�.�0�v��x��=���V֣��zkL��=��ъ:�W����D�&�S,��4Do��Fz��n�r�	�ӡ^�ae�63��qyH+�~�$!��9��j2&|��-%�x�So��J���v��,���*��s�� ��T��w�)>Յ�9��#:��a�fS�j���:�S����7ɎH�ڡun{�����R��`��7<��d�R^u�����9����~��P��\NY���M<,��l �%4�#1�5���L�=��>,�T��+�[݆���<�{(&�^.=�+1����s�ݨ�*)���;ߚ��T���q�R��!c�rI���I�<ϟo߈-
��,��	��"v��j
!u���!��n&��<��/�W��>�څ�PK(yY?�p�v98K��s:��Tc0vI� �(�0�ô���o�P������m�+����/5�Ա�>c�^���������&������\o���d�|kQ^d.Z�X����}�u!�2�؀�,��܉�Z ��V��=�/R|��F��hc��R��d��Ѭ��Ng�!�Jj3��[�%vp�Q7\�A1��9�������W�K����f�uF%e�.*�$�����I�\*)Yeٔh.7K���(dGM�ΜK��)�\K;�â�0��ץ�e\��Y�xK�]���;�e���q����%�x4Vm F��n����/��$T�w/��1����r� ��"*��i�\*���#3��)�^8�J�F������G�_�l�:%��hE� ��&R
ȥ��~Z�P���f�Y��S�%גU*#ZW�9]T*�5m
c�����2����˖�Gvg�y+adL�e׏��T��2"��g�$J�~���1<�q���A1]Dep�j��"L�J����}�t&6�Z�<�}���H��.��~�n���#�;�eP�����+�u��#p�&����3�_���r�}�M1E���6"����c����Dy���YX��2�G�W����R�(/�?���0��j��Fwp��.�����n�������ƈ]�('��8޶%�h,��$�>�a1�c���E�_�-H�/T�,��Z�Zp7�.��nPW�BZȐ}��Sp��]g�h���1f�lCm���ѯ�<����Z���!��3JGz�Z.g�D6IX��o/��/��kf.���^�q�C���g�E�%u�g��);eNx�>�E�̠�������[��$8����!fĪ�l�u�zDt���VMqbYX(Z���Ä ?�%�r��}��CT
��Ɣ_Pv-O���|�i;5��პ��:ūJ������r_o��-;���.�؏�h_��xI�c ��ٚ�;_[�<��b��ݲ�"VyCz��5ake|~����p0{�O;��&�(/�g8��'����O����U麐�r�V^e71����w�jI6��Z������}U9���i�7�t�=���H��`�l�\�}ww�Z�I�'`�x�o'�٨�.q��#�;�q��#ŶO1�h�~yd�*m��Q?�6�5�i��u�:k���q��S�ѿt0'��A��i50_��J4�T�LݹshuWMpn����F�(�?����0����GC=sઃw�a����@�h{���k	/�tE��[V�P��Q����0��\e{����t^�e�Ѧ�p�R�\z\vo��� 1@p�n$���x\����e�˻��l Ā����A�i��D2J��]��#�} ��+ϥ�Vv��h-YSTI�h]���e;;����ߤ���.�9�ת����T��H����@�(�A���,= ������>�`:�5�9'/��J����y�sg�0w�586�g0�@�u3�'�t�����DO���Hk��kw7�� ���?YG���(�ue�P�Î5ߨS/��Q�1��e���]�-���%��`���j��Mc�f�s������.��*Z#��9�����֑ ��xvz]�i���)��[������h�S�+x�w���&}[�T��0�!дylurH)��"6/��A�U0��/�W���[�)�,��H {o�e���q� h'���1$AV����V	O��C�H� ��Σ����]@9V��g}�Y��x{鱭i�(��I�-���X�x��~�5-,��)�V�"���5�a�ZFj^�}�)Q��e@e�*�5׏�q^k"Rp{^[g���x� 3�ο&�������M�o�*��:��p��^�t����\lj�w黍۵����g��z����Gbp����H.Յ�l֥�K�4*g����yuQ%Q;H�y{�FA�K�T)��.�7�k�g�|[<�/+���;\	5�)"i��.Ԣ��L�p23��|�ǃ��콸S�����ގ�Rj�e����\ʦ���>��
S�|�&t-�^��aIbY�+_���	6fh��u�h�ˈi��~�\�E�5�V�.g(��)�������GcaO�^a�g��1�t�����F%��κCP�\O�?{��&o3Z(�w���e*�H��Au"�c�<�T<Z���%w+�3�?���MJ�6%��]���\�x�����i]-9�{�{z/�w-��S��؈p/�dM��/�h����uV���e�����@�[R����.��2m_V�������.=
B�oe�'�p�������(<��u����o��	�Lq�f}s�p�Cr�}`�f_�,V�$\�|��@����f6N�.�s�d�=�u��֠����s�N��ĵ1��Z���p��ý�6�X������TEu8��?�;X� ������U�7^����luU�B<@�lS��l�@p�k�/8�6S>�ٲˬ��u�{�{a�n{_�ڢ>��Z!v>ؓOqݾ^��K;>&�#z�	�J`~Ȣ�pVf�/�}f��f��$
����(�/47N}���,��=�nR[7}� P-�u|v~�����1Si�Y���=R�����͌3�g���5�U���8�����E���g�(��M� 0��+7�i���_^���s���]��᪼-�D!W��3����<*%b�����F#�,�Qp�P�'���eO�8.�����cjs�Km�eώ�/�=���4��ma�qN���Tkv�X�x?^ڟ�fe�(�!����*��FvrgCIġ�%�u����%�((���5V&_m��)�4+�SArx�����L�\��N�ѷ�d斍�b���y��<�[O��a�yU-�+COr��� 6<ݮ<@�tSLY9�+vĞ)]}�+@��"t�ӿ�rԣx*��2�\İ?��_ES�v?�e���Y������L˖.��IYi7N�G�B��\6���po��Wtg=ö��D!偖�T�A��o�t�$v����`� �O3���V�<rn<U���UJ�џ�?�}C�7��D	��ҨU2&�p�*ؕJW��2�*�g�ϕnO��
0��Ǝ�9�#�k�n�0���_m��p�OcG��<��	��3c;�)ߨ?��>j�����C�5�|��[��6|A���N�@.�D|ń��o<��V��X��/~�,%�p����b�j}n����F�N�e����i��B�xsX|ր�f�2�@�މ׼��H���-����Gx�۱�2�h�����t��ݲ,d���������ٍ��[����"����%a��`H8��]��ء#��@��Ȯ5��y�bF~�z|��f�ö�|��g���N��B��'?l[YU,�-k]���޲�{�>"=�i/�X��\y<���1��rt����tEF��tU����j��̫w��KC=�>#|W�Y�� �e�j��\JZ�O[ȕ�'�Tg���{q:M��975���B��8\^��-O{��wp@�|��Y���<��L�c�7��t�g��Զ?e��2���(�:'ѣ�?�Ԛ��ћ�v�y�ԛ�g���c��P������_��9pht@%R��~/��XK������aB=?��`�M̘��p��������1� �1L��$#��B��:T5��~\��G�F*�E���7���s �:/m���{�|dM�P��&��YhЎje�$y�&g��)���@8)�����bmQA�7j}�9�ǤZ,E�(�pkh��VHQ�Pk$���zJǕVn"�Uly�� L��gϴ�o{���43l�r�C*��4��4_���Pq�:%��PJI��7y�.�NucV/j�Q�g<�ft��MML$�i	�N�$���`��d��5��}�.���p�i}�-!Q��t a@sG�nSV��&�E��m���Ty�&�Z��ZWH�_r�����L��q@�U����b�6��6a��\HHT|aƪN�YƇ�8��'Ǆ
������mƲИ�_��2��Ekq\k��:���l������M��� �����Ч��!�Րύ���d����*��6���������o��|�>��S >�^��:�S�*2��{�ds#���"��7CL��ݒR��uS`b�xX�������c�)���e1N�!�9l|��g.SM�2����(��D)��>�O��`3�-Gl�=��K1Z͑?oDf?Q�I)�OL�c1��g��'[�< QAT��l�R�2`B������Y��0�˔#��m�� K�Ailb�{��}R�&!�b��vmPt�c���@	u0K��Ȝ/G٥��xK�:���!\Ut���x��Rn��ze�/8$��e�Oك�LsKl[��H����[2��G�x�Ҏ���aG��B;�&/���D�����W�wB,߮6>�5��r��!��~;�ۘ$]��������I�[J��"݅Gk�;¦\�K$��Sve�M��مuܙ��.p�e�A�a�m����8�QI���z��Zw�cI���M��Y6�;�����f�z�n`���筝�V��������o��.�TD �=�V�t�������;l�.>Ԡ�!��Xu�S���[�V�Yй$.V��G63�~�L�k5��ǭ�ȥ�����2���v	�/<��R&\k���	/_=K�gc~��H��/^(���G�׶�M�+_�ͰU��&��='f���.�HMK8aeC�-��t`9��r�t�c�c��������H�����2BEE��\ΘUq�H#���qEeBMyQ�Q�B^���u2�l�D*%f[���e�W�ė[����ބ��w�^ ������� �Qؽ\�yIOxY��W�@P �H�8�q�;�3��G�7���*=�5	@�l�Pg4����8ރ�d1e�IIM��zs=K�h��!0޻��P��x���4���+D=��=�G0c��4�r֭���3ml/����i���㯹n��n ~�1uݡS-OQe1MS/��Q���s1΀1�5�9���!� C�9V�Jh���G?G'��BR0;{�B�����Yp��n�c�%Bl���$��ᣤ���	< ��ܻ'�[�`�o} L$�hk|rHt�����=I-��\�~E�S��l�ߞ��@){vm�y�F�U�6��@�W��ɇ��պ��"	/ 8895�i&��S`HD��v������@��T�
�Ƴ�{�:��khi�1Ӽ��|����>\T��,�z�䮅)<�Q�@�@W���k���ܭ��z��n^�o��C`{*���xS,��軑��Z�a}�����P`V���µj�Jb�:V���	���;�(z
���`�[0~(�.��`�eQ}W^�X��kp=�'<��>i��_�rL�J���(�0�?���*^����\��b�`�/,�=����os��"<D�ތ癣ݭ����Z��Q��`�2�}mu5�a��P�X�	��RV��
i�ͪ6:|���8��1�Q2V��QW�'Mɼ��r�Z�OZ)=s�W��R��#h@�m:ѫ��j���<�� z�A/[����<����믅--�i�!��hvRRrb���K�M�.�T��� +�7��A���������q`-���)�n��*+�=r�m��꟪U1��i��hw���7�U���a;!1��'DO���E��*o�B�RT��������̏ �(����d�H�K.�ߖ��O.,��8ߎ��U�W2V933�	�	�-6���ϓ�)��(�kߔ/�n�ųHSgI{�ǉ�������˃//p��(^O�`m�t�ɿ�|��ΰ5���傔��3&G�_�E�\�G]<�}�=l3���>h�zF�����_�ȥG=�D=Ѽ�IF:��ຏ�i�UdJ%xz��W�����9�Dv���t��в'ɒ�����7�=��j�|T�op�D/�"���)q��-t�{Upѫ��;#��q�삑���RA�Hhr/|� ���`џ�7`�,�.���WJ���`�υR��;r������Q�����AXm�\�b0�S0������9��a���b^
%��."�:��	��r�C�	rD���ꝸ<����#�Ǯ��fGzerEOF�v(�$Œ��U��f_�q��sB�u�-�.O��/&?8:��E��BMIX��H'�e�|�]����Ħ�/H�S�٧��V�l�/��y5�sq��j�he��݌/��y��Iӕeo� ����1���gk[F���c���q�2��9��K�̅4N�ݭ�ƪ,�M�.�M��b5��/%A�y,��wGV�{,�GКD��-�&-M�.��n<��hv2��\|XX��Z�A����9-bxxx	<E\5� �ڲ�OD�^ť'��Ȧ���"p��x[�[���˲ӭz�C܃:�ٵHх��^�<���0+�56�E/�D��Ũ��8���*`0 ��̃i���ϰ���bb�+&�:�Y�U���LMMkڙ
E_��'�Ƿ�0���Ɣj��W#|����(�
N��A�=-�e�A��>>=�N>0>���H����v�V��	��0Z�$*�|��f�ZYY!N��w�	u�X�."|%�YZG5�F�hG>-T�Q��uwu��V�}�J���;���م߼�h����өY�9�*='?�V��%P(T�ULJ
<P�:11�[�_���?��0^��>�k��6RY��	���y��y��G�x������u$�7��kqU�p�ş0J�2<�^�nh�	;zӐ���=�n����.P��TǷoy���7!����d�k�]g�`��B��d���Z�qh��X^�� ��'�b1Ñ��a|$��lCԝԟ�OM�?;�\1_�b���j^7jd�N�y �-���x�A��M�d�zhϡ�9Ɵ��ADh�k�CZ�hj�v�Z��χ��q�=
,����������L�2˃XyM�8(G �eB�ج�o|��8謼���w�kz�����[7-�3�%�r�s�l�KP��_m6�ub>o7�
��#�Z�7hU��<�'D*R��]ID-����]��B�6%	�iw��}۲��� nn�&����f��D�������e�\j�ty��[�Φ)�ܪ�:�,�}��L�P����zY�c�ɥ.z�P�H�����x�#�������}=-44>��_FDn�6N��ʹ8Vv���� V8,��H��J.� ���|�g�5ӬH���mJ�WX�}��6̸�aFk��}�o��FE���H�B��Qsp�[��h[���e<骎!!�%��v���n�g�qjמ���/|� 'i�#��8��nG�`S[/]�E�$��']^��Lzw˥���z!ºa2W!;����~G��O=�����?}@��	Y�27\<�%¢Rv���e0�9��B�]��\����.ZLwE�c�D'��B�8F�}��{�F��g��Jey��Y����l��}GV��uq�'�G����PݕOW��:����G����R��T��=��kG�$�&&JZ{.v*${�{I��S�ӄ2'/�NWRSJ��;�A�g���ݨ-�����y�y���g���
%��R�@����U��z�f�9�����#j:����e㌲������9>i���7�z�=���_��p毒E������f�T��w���a�G5������CN��D=�����g����f���_��}yX���1!�95�3o���_�b'<MWfh'��-�y/�ԴC����af��s���R���>׫�x;�>(,�u7<P�д�1��[:!!�݉苎��/��۪��4mu��l�I���)�}xϤ�۸�.��d�Yt���td`#W���Q*k��X"�`�J������M�d*#uK>����rb�3&* ���)v(���fW�݆�����=WiIt��w18� �`OS�J(V����$�,11Q� �����&�fACv�|���p����l�~��Q��@C#����s64�Pr�������{l�s˔[ �����ZxΈ��L�ݦ�$��h������|g��ǒ��@:q�����n������}��#����=�UV�� ���Y󈉿J��8���$�����4�H�	�hD��v
�/�^;\ }X��N����\7�z�����<P��`���Y�
���iH�98��[O�ݾo;1��	\)Ml	��sp�[Òz�\�'Xt��#җ%S�b����6f�>��uu�tŦ�ݶ����mW{qo=�༴��2h�׷<��&�S�;:4eh	1�*ߪ﹌��\��lͺ��)z��0�w;�Vm$ ���Q3�p�ƥ��o�1����9�����K�c����Q�v��2%Ie�tl7���\���B7 ��a�?�!�a������ٖ�P��8����|�
���1=ey��#�%��O�p���)^f�+L�
��t��.�� ���
p].�L��f�{0�ż��@[�`���(DN%'>�;ʵ�?��.���LBЄ�����C|�t� ���H8���-l���x�B���s����>�)CS�O��#P�y䢧ݨɻ�'"��3��� $�|MHXrn��ˢw\��!Q�=2E��7%e�z�q�jr~�g��.���a�����Z����>���:D옟@_�n`OJO��z��	eD��A6�9�*C1�o���G��W��3�w������U�G�^���)f⤭�<�\xǦ�[��B��^pD����7�k�!b�/KA�_�^m��1y~x���KF�-�g��ٍ��������Є���I$Ȩ��P+�q��S��D�m���h�Ք�@ ��\��{0�Ii�Y)��sTx<�l�A��DS�g�}�o��~~hHy����/�(N�0��x�0�O{���9���@&s��i�H��I���)b#3�M�/�����w�}�D5�8k��z����u=%�u;��o}��%vrŢk��7/������_�y���Jּ�b���(.4���l�(��U���6�~��4�'�E�|}���d|��X�R7��lD�׊�nO�ybY���vBd'��mB�@ߔ"V�-sel�Zk*S[��h.IG���ąc�KT3ڴ�Q��jWrB4�c5*�N���o��I�D�>��״�?\����V���
�h�M�r�)�8����Ѣ��Ngۘ�$��$�PK�n?���C}��7@�^XL���
�=_�Zp��P�hA#N3��@<���9E{#C��I�"����v8���9�UD��<j�EeX��=����yl��L�~�z�7ڬ@���A����4�i7;�6VO?��7P=�� ��zB���5�m՘g�)M���|�l�շ��L 2������ax�V����>��>}J~�/��J"��#/"_[���@�� ~�rk��K���i���iưe:��?��X�`T)���Hm���s��; �k���!Oc(�����zb���+ybl�?��'4:tc(�s?��ٚ�|��cv���H�~������\�kg��Mڮ3	��>Ҿ�~��kKI�E��.�M��@Ko�e{�Jj2� �վ0�P�?Sd�+[FS�͡ՙu�a�!?���7(Ȓ8������K��x[^��o�o=u]?R�������V����U+�a��3�gJ��D�]5��GS3jF7�`lf���uH�Q���K*x�
C~]O�܅]�z��F�kp�ff�?�b�F��
� 7E|�7��1�@�	�C՚�q2vU�F���<�U�t���a��Ǆ��s����2ɀ����2��7��]�!�+o����S㍉� �''�<��k�_��U�%�`~��cgSŗG�0�/�u�t�3p��49m㊿"T�9����2�q��Κ�}��T���e�C��N�Qr6�nM��<w��eLp��z��
��I���{8��l}z ���3	�n�(�1@���3�u�[s�~I���􌱦�)�L�����@��ܴ�|�Y{��|}}�����5d3K�u�7�����/G1��5��@��_��5���^ღ�W��+C���Su�Zz;9n}y����:�W����8C��;�n�?�u����������d_G���Y��������w�k�w��V���wH�Y�Z�#g��;�*�L ߣ^����l�O�D4ey٩߉D�����В��%[��BsV�뚬 �q'��C�(��_����g�bʟO�q(�^okl��C>��4ט��x1l��^7u�vwݤ�C�;�Y����I���p/��4�@T1·]]��}6P��[�1�z�ű6}gT��Br���j=}�B���M�Ok>�_<���O���%%%)��LE��7�G����ݺ�ļV"�y�O����6wv���-�m��hXk-M�B�������ML��Jl��$v��<;F���Ӈ�,��bs��}�D6?*я�jI��Ե�RYI�/��� ���u���d��xe�X��e�;Q0������-�^	E���;���:���5��ıWYf�J]�M9V�\L�L%�������?Z^�O�_�q��ʗ
n�\V�������s��]W��.�ض�i���8�N�9m�>�������I ��Q(�x�y�s��t>���t����K��� S+x8x���u���o������X;E��1����h�Y�$�ϭ];��>�	@�C����EӺ�֙wh���.�]���T��B�V�H�i�����H��wO�ۗ� x� ���n���w�&�<y!��c��)Z��x�q �S�x�2��_u�-��iwX���27H��$ ���\q%�U�xۑV���8�t�%�10�E*Đ1����J�6G㵤gn���6��B����� >�=;�
�N�)�Fه[p��!�V��V�tL�{�kGW�/f��{rc+°�C'++Y�`� �8�����?�Fp�)�d��#,f����������8IKK�ى�

�f��9�+�G6���4`����Ht`
��d�Ϛ����E	JJ֚�����Tz�6�Ԓ:L�����{ ts����=[t��{�U11�D;��J-�C��t�!'�}n=G��)ˋt�㶑�8�:�S���^w�\;\{���V(z5�
=�@�\�#e� 47�C�Rb$� rc�7g����F�ͦt8fN��u_>�"��yQp�x��Ծ�mӖY"Yg$���n�\�<�'*Z������P"�`N�,��F穲��5��#ז�����D�kh��WoW��몖����o3pi���M�?^�W�08O C�ı�ݵ�q��췇�M^�;f���{���d���a]nݧv�^b��o��UF��BEGI)���b���4� ϰkS��ݲ߃G%*U�G�
��Tj5�t��zJ�ޔ���z�$~zL� v� 55j@�4�t75�^?�9ܲ�j�.��ދ���0e8�K8�p���%�;~N�p��Uw5���r��p�ȿ�|{��\JUT��5�K�Ąu��wBC�^g����fU���.R�i�_�N�^4��O������͗��k�l�Sq�V����i[�_�7z������z���w*���+MdG�gO_u�b%�<�꺱N��F�螣G�@P i+��@I�1%y�=H�������Z�7�2L�.��2��g���n�T=,t�-!f?)3�uY�t�R�9���ԝ۞��8 �a%@B]Nc����h
�g`���J;�Qnnl���/T�&��4�e|�;�+��2A�w|�q���i�Y-+-� hkر[z�:��I�9LU맔κuh�\�Y
��t�����V�E���>Mڟ�y*�^�/�h��׼�p�}�ۀ����ŵ������ͻ]��������R�?)(�����+2I���O- z�(���iMXZz}]�����~š���&4�H\0��CUM[�C[�����=�`�/i������������2�_��Z���7�7qڧBi�ox�O/1����>�uW����wo�il�}J�X�{y5X��M1��������~[��d��MIOQ�ǥ%�L�Ώ�ф|? \�"��qV`c��OVC	�sQ�ǗkQ�;q �Ŏ1_�[�:�GNn��ϟ�3����$ Q�s�?`E%�)൮#��MRw>K�Ի�K����5U�!�OK�J#�Ȫ+�a��Q��#� �w��m��+���/oX*��2
��O�.}
qt��L���\�E���X`�o�i��������QQ�_��H���� �݈ H7H�tw�4�-=H��R�]24Hw�=�����X��5Xp���|���{i�;���c�.��n���,Ro�J�fk-��J�m_G�8P:�+�k��0
��z�D���cn	�z[q`ٽ��tH�����ڔ��/t�{0�,�=�Ck ��n�H>������:��ѻ��w��7ʪ��'����h���e7�tyqO�C׼p]�v2��R�y����������511����$�ˈ�i���ƻw���,�|��,<=S�I�|�������N���3Hm��6���}i� ������G�W=$\2$x�#��J`{��N:ۃgX�>��HY�׀ԟh��WYë�hP���j�!��<�m}ML�e��gy���*�z�]�;O�M�!Ȫ���Ի�yf�l�	���,��9]s��ۓ�X�-�Ow�jV����}�y�U��D0Qe���8n܊L�\~C���?� v������6"�	pa���������?�3���X8�O$R!E���V%M��;3�7�_�k%�p�.�﫯�K�'ةUe���~��q���b�z7X�J�VU9~>��x<�\��\�L�ч
��h�ri@����a������pY������ZU�0��sK�A�=�����Ő�H T��! ����� *�-����OOmmЯ�ƺ�Sv����V��|�����uR�k���m�4�b�!9EDY���J�(�z���S3@1�lK��E9.�����];[69�����p��Bm�����r���Ђ~f��;%\��Es�OF�A�����b�,SL�i=�i���eqs_���(��g���(���Fb��3�=X��O�LYC!���lOP��Z��83��l�2�8Q:i4���2����<a��VO���.����&+���"s�N\
UG�S��݋wR�m����㬭jj�y����+���\�*�Se]��A/H�r������ĺG�B	d�A8��c21YGxn����P��Sl#�px��5�/8�ٔk;TH����������]��:��Ǜ¤�16ğ��4��W���E��vaT���B���j��H�>����=|��jjv���#I��Q+�n\�j�TWm�4J�+���?U1lL�d��.? ��j���	��o1%0^e�u�����o�>��b�H.�ߓ��=�6N�� � �Ι�ݯY��Ϯ��q�ekN3*��a1_��KMÃ��LS���*��dBv��p�n'������5��`�2_����B�[��y�ns���v���ߢV���e�D���~�����&����d����>y���q�� 1�g��ƸV��tQV���:����n�Z$s�s�k.gb�^�[�h�5���f�n��o�W�)�:D�T�o��l{��n\�z�&�眪��Sĺϱ��3���s3w��㚿�%4g��]�=X����|�t�j��5��`�PQ�͉�Ԃ��Z�¡�b'+NΟ[��uC��'r�c*l�		��M����
)�����J����US�	�dZs�c��^<��c~gyh:K�J52��dԐ�д�����V�pv	$bpP��� ��pƗ2l\Q�����+�L3 ~RǏ��h��t4��Ŧ]O�lQAC�,�16U����K"�?�ų�yb�۾�n����YD�6Ɖ���;���A<�_4�J�2����O�]���-X���c��R�Z��/R�Az��lߌ3��������4B<��3�;}��4R���T�ux��5�"�'*#^O�g�7B��׆�/z�>�������@4�p�@~�8l�L�)2�q�DE�Ţ��'ϡW��U�|F�UQ�oP���ob�S���c]���ը��m�X\��Ax���'�?*��f{>�\��;�t��Yƾ�����$����!��]1P��3l�Bz�&$$?�ۙ�}U�$Ϝ�r�r_Ub�C6�'"eS��T�T�id+���w//���_zm������/��Z���v�j/��Ч�C�(5�5��yƦ��UoN�5Ky�]5n.N�mOw	�������6Aq���s����
�mE��5��G�>e\���Y	Fe	�w�%��`�����7��iD�|�\���>����*�A
��-���G��O��B ��@W���9�o�'t<;�E�:I���q^�4�.����w�1bQ��9
� SX��{�/�F�s�"�&��������qr]�+Wttt;oN�N�ZX�8e��C�ɨ+F�w�f�0�qk�Ӳ�1f��^��e�% ���WK����o����F���	� �9QҩS��9�;o!ӿh'\<�$j���ג�:;��5�>��_��s?���̆#���ߠ����G����"Shf0�ve�^���S�Y+�*4s=�0{B��dD��_�(�T4�PĐ�YurJJ�����BLL�
n���
&h��.F���rIF�jt��=�C�ʾ4��:����Ҥ���C��ސ��;'�c�p��]��R"RR߾�!�j��	���Y푩u�X�G{����{�,J���hk���.���������8��֖o��\��
��+������QZrϣm�^<?l'�0��Q���n%s��!"W�"��M����Gc��Y���{WBֽ�&
0�J��ތH�2\��`�X��n�[ėR"��|Q �P�H(��7ˢ2D^T�\W3��/�}����-)r5��2>~	s[�Xӿ31����p����z��>(����6����v-5�tA�V��G��("a�G���t�G�K	g��%$��E��=K@��{���TTt�+��!�VFg��1>;�.N
E�T
�K7�=��q&b
�l�u�"��}��>#{�<Z57!����н���t�Jw��ۖ������U�'n�il�ET�� �������Ky��~^�����ϒd>x"w�1�n�z;s�� V��"��"�5�J��i(�q�ˁE���/�Q���K�_��K*(`�2�44�#{��w�����u��S��_�vz��ccc2w��b��a���"��I����/&=��'�5�]���:���
VJ�o�"�Wn.�/:Dn:L��+?kNp9"gH	;�!��)+�)�2��w}�I~fS�թ�A�����s~�ޙ���J��#����FB�OE�����9�_8K�^�9�޳���\z��sً�&X��ћ`	@"��������Y��#��
���[9q��&�u�Rd�_'M��c�;��4ajj
{|��ѡ�h�Kc�ڀ<Gv�.�Z�>v!��B���|xl�ӑ�l�".���	�t�%S�;eJ���ĜI���NQ��K�+�ٮ�z'ۤ���o��)�}�/:c�U��ĄC����uCƻXt��"�y=�w_ J����v}���~����Z/�AdNgˑ�[K[,'ҏ�w��~���\�� ��C�6�7����^���M��ԡ���iHL�b,�\I����K̟�q�"ݮ�7��=�b�v�D�0 �GҎ.��V\_�{�͘U���R� >?���$Q<�<�G�7��8l����ˋ��\�>��Ҏ�+��y��)<�H
�:\}��F*ɹ���uJ3F��9v���F�֪~~��s��g����C�:\���>JK)4����q0<:�n�eʀ���L�#��j�A��E�B��L�mR1�a�S�wT��{����ɚ��Z}�z�@��c�X�pJ�V��ML���r�VDU�.)i�h������^�������׭O����B���\��1"��R$N�J_���ȊEGw�_M	�u�ϛGh��.��E�b"ަ�;�y*���"]��!��ၛ����ʈ�O������;���6i����OTp���@��5��y���N��?ے��k�	�)N;;y��D�,�5z;��^U��N��_�M�Et����q��i��|��e?5LEN�c.��_fF�5
i�0e,��)��BTD$C]�a�l:x�ͧ
3�X.k�#��	,���D�c�첅'������"�Ps��{�}�ފ�nӋ	#A�5�Q�m⓬�3�D�i��J� �!�G�w����6��x����|��^9�h�~.�=�������KӏÛ���2����Dz��w�r����Gk�G� �����0&���+�0��.�l���I��s�FNV1����`U��h�����p��M�B����@���V΋���f|f�o���?Ǆ.γ�n��2�y��OuU�ڳ}&ː3d�E`	}^��ó�}r�>N'�7؍���x��]�l�}@��7��I�lez��i�f:\ѯNk|8�O&%]�PL%�$��Nj���®F��
�w��.�~ɉ6+�����\1f�c��]��\+�˰`����l�̢7c(A�4^��n�i�~=�01I:5Xe�$�ڦR��~�C��݊%n�d$�ٸ$c����U�.����o���Om�0y��~�Y[�ȋp�4B��a?��Y�?�z��~�n��?�}���弯/�60F�sI�O���E���/~��o�{	��`ϻ���^�ę5�@����	Cb���CE�]?>E=d��c\P�hr^��������/�b6,W+0_
_��{��'�<�e����U�?�mʦc�/��9�p���uzk�˥�2�«�����*���"�qY���Ƚ(�+g{��6�ܿW�9>"�5��+d���~zU�'�#4TȆ�\$|<��G�M��|g�P�����2��czD~���1�W�(���]�����3�J`m���2D�����S�scp�D��2�& ڡ���k��������
�E.zx����s�5s�f����v-'���W�c�g�-���v��a�A
ގ�w���kA�
5��Dl��7W��w筧'��7w��V��=>����{��#n0-z���[|x��𘅸��\���c��ӋlE��-|9,!��G�
�X��+Gهm��\)9�>��@��z��Z�6��H}U�o��_DtR2�9�^*Ȯ�g�Ǽ�@a�\��z���#�c:����A��N��� W��h�)�����r�h�RS+_��U�Uj��:2j�d�/��4��a3����:l>q����
xB�G׏/�c �_�ίs,&�VX1���f�	Rd����5���;ׄ�q*/G����Z���h�B�l6, ��'�5�H|D�U���R{����5Ƞ�����u6�qC�Ƽ�窢���������+�q4g����(�Vjb���5��ev����?4�:A:G���悼	�����w.���棍T�~���q��1~\"2R �/�~�5�Ԝ0lz�y��G� m��K�i� w�K��^.�AJx��#Q��]��'��%�+צ1?CbE4wx}+�&>��HQ�-��o�89#�sgǺ3WD�#B���U/�SY*B��-�*���!B�}�:ZC��%*�W)*��z����䴴^m9c鋝���:����A|�n\8]�7��qZٳ��_؋̏h�T�%& �E�rp7�(�"X�1>�*�Z$��R���#YɨB�ƥ�)��c+�tZ����_5^;����f6k�����܌��H��>�^�::k������'ZkST̖�	t���<�hqb8@WW5�d!K���lH� �7-��r���'T��z�����r+9M0~)�
:h�>[�G������{�J���TIWW������2\$-����B˯�ηߞ�/�6�%��󅉡�ll.��p��׏s�˱���.'���m����#��'��A�HY,���.�]�P��Ȟ�0)nlF��ٓZ|7�l���#h�t��uk^��aP���)\z��XO��,����yv��׫~�Z�h�H�����v]�F\>�嶛�b>^�zj�����A_"3��"��`|lj�'��@\�x'mK
��a�o����Tgg2+�@6������1��łW��5w�XЋ�X�Mܤ.xT`��l:r�utE���v[+���[�{c�uo���������KՌ�׏U�ʦ(RR-���X���d��_C�'ss����>�,׷D��bff4�_��"���l�oT��eoi5�����&�]�����6F�&��C8��(�D�S~r$	���������]�A/��X����G�zu����D�2R��J�c��kw5iԀ��h�j5��W�o0}�ND�ד���U�������W�̇i2Bw"w]�PH��B`c�MU7Y��4� E2TI##���+�7VO���X�:u�)h=����鮪������2�/5}c��*;�X5��ev��as��/-P�ְ��5�����;侓i[$c\�urv�\�פ����2޻��As��{���9	� 0r;���:���D����iY?~�w Ʀ�N�¢�u�<�j�H�'�lCՖ�����g��|��ࠧ�?4	%VVV{9�����L&%r�e�8��H#�v��R�-�S���g��d38��ߖ��8qCmS
�ݥܔi�1{xYY�g�dM�����s�J������(�Q�����z=V
�"�ok}�[!��_C������t|y���3��N�b��"�adg*��.֦���궻�'D鑹�=e��D8�^��状������_S�;��e	�wգ�H�}Yi��@�6�<�������*�./��6 ^־�Pe�Ƙ����At�S?� ��7���*�!�y5=[�F�\T_?l�a�QJ��
#6�����pu]t�/��)��(�1hZ*�sg�˩@SM���S�yjH@ \: V�INcg��_ޯ}�%~.'��x���v1�_�f���.|�פ]�lw�.��>�����?�H�W=�����X���~%�Y��W�gb6e+'J��P]天{)۾������#\3]h?b���K/�X�5�l������Lu#:�H�:��W��ل��m�����Ϣ��k���﷪Dx8g7�O��x�
7'�3�:W��`JD�dݕ�(0f�F�f�����hc7��G"9ش�JW���?��#���?3Q��ظt|	��{���a��#��H� QfF:�w6���o��6Z�rE�*P|�o� 3iLn>ЖF1���%1@tF_�RƓ��?й������'9qY�@�(<��:�����=��9�غQν�ڛ��5Zy� ^�`���_�b��v-�������W�j�ou�2�q��hf�s(����p��ʫ����}��h֧�f�zkgǂ'���I,�vv��w���x۝��Ү_ ���Ct���`�/>|�^��	�Wo߾@e)S$|�U��|��Ƴ�gE �[��5�/7f�;5����&!!�k7v��d���":#@�2B@�P��i��!�]WJoػ���9�%'Һ}��42��k�4;Q�6AJ�H��򾖩]6�RT/�]Hj�BAIU	�r�A�@�N��(Sd������P�]]�k2~�3���_��L-x����`5��q~���h���F����b��<���gg��aj}��"�B�M�ڂכm�2	Ȍ� �"O�m�M0�	�R>G5�.��z�w�L0<)=�䯨!�}����Ԍ��Ы��E������81�8��p�t� ���Zy�x0��w�8�Ԙ�qqh�g��M��]�K?�ڔ��V���5����|����{MM�Yfy�sx R}pN��Ki�|�ϖy�[�qjjj�?F� ��I�õ��6�G��]}{�)�?�����ʿ�"D�Z^����[�e`��l(#:j��1�ȼ��ڭ�+M#�/�ܹ���坑<����%�u���s��MHϐk���^ �K����禷4"kR"ᚅ~PG5�|q�ٵ:��h؁Kn�x`��׍&Y�9�L�'g_CH�:5L�4��2�e�xz�\�1��TX_�	wN�Ӎ���ߌ�E�t$�;��@ԡ�r-/��^�ϸ���z�8Y����T��5����{��e��ܭ ��F;;�-dK�V�̚�(��-�A�Vu?�
[a5c��fh�0��Fq��(���0�y/�_b�8%���~c)��E�]_q���g�}i/�l�y�$��� �ky�7�5�:j��k�!��"�H�הo]7˃)Ajc�'2%�Ǔ�3������+�1DE�|6���㚅&4Y;2�'�!�$�Z��0~r]�]�kDRΤ
��v�t��G�z"��<;9Ǧ��=2@���Ҵ���jE�KPH��6�K�uTw��D��%F[gR���%5���fa��~`G�=��r�����="Y<dھ��kV��Q�{�4}�r��"ML�����ҏ��pF_=�.0#��5Z]|E�� %?�c�1�����=�6T���]E]1��M�`h�)��t����;l��ݳ�4k�����0;&�w���Q�d����7-�[zܜs�3�1��MO$��<L�r1c��T�\u}�@����,��U{bgܹz(�\a����a"Z�s]����dh�b��[q`���X��W8�u���Ӈ~��Xx��Ժ��A�%t	��(�9�\��8��ޔ`�Z�D�a X���w+��""��G O/�JTJz�J��p_7HЋyבb���(���c���۽�cX?�Ci�ٳ��A�}7�oL���C�}﮲���',B���-�,���������'
.��a�J�[�-4�d����aA$54Ԩ�\�B�8He��tb����kr��U�;x�K�y4�}��e�Z�xy9l��!?$�t�$�$=Z��d��_۱j�c.n��0l�{B�����PR����B8����-w��C�c�w�?|�6It�\�n���#���:���|��(�3�b�Ю��wY[rսYUWR[��A�vu'�_M5-�|�;�gh�?�����yuf7Đ<!��0_�Ȟ[t�g�w�q�vrZ��#��!Q��m�YO~����ֱU��5{&��!������+�(#xA�Mw���8Q��`#�{8۔7�:�HR������Uｆ~�!�߸��w�e~����	�T{8ʗ�/�ł�x3�Vt�Nmi���ô���$$�(��/ϰ~Rǅ���/l%�F�|�T��tk��\�D_𘛳���c1��Z^hh��e�;/��H��j�����܏�֕�s��wW���w�[o2�K�ھ��tҎ�L�9�ϖi秋��{�����K-n��y�L���d�8��[���v������9��þ��!�c��*zI�Ym�nw�J�tuZ�?Er��~g�2�L���>�`��{����1[��0d�n�ϗ�W_y�Z��SE!�o���v�yTz$�?M�N�hV�$���U����8�-�������y�}�Dj�Rh�.����%���N}3�c~'�wr�8��2mY����������濲��O�J����^�6�*�>품�=��(����z���L� I��	���`dܣ��f��w�*���,�.o!6�(� w���;�f�r>>~�w����Ǜ�u:�P������pwe/�����_�䛱,�,��5��j��ɺ��x�pa_����T�$�1w���]���e�tr��U(��3vJ�&-Gę��� W��}�sњEV�5�p�i^��5��hnqm��l�K���ϧa3��{�lpim��l��LA	�H���v��jԿ^�DL�Ǝ�̰�b,е$��j8-��T݂�g����@J�%]����qMJ��;�/�{�2���H@�������C\�m�{�?\�G��P�B�}�_e��w8.�e�7~��`b@�4���o���P�}�i���XѬ�^w�}�j��L+��o^�\�
�G�s���(��H��퀐l>(L���Uw24������b��tĽ��K�_taPy���جLe	���b_s��?�a�߱'޿?��K�oЍx=��Kv�Ɓ��4��P�L﾿"�a�$�1X��^��M��Q^u�bVFS��t��n��1�[�vU��Κ�{,��=��yq������Ⴂ�|��	�5k�I���&3�4��~>��|]B`�l���8zS��j�����R,�Q �5�̧�B`����am2$q7��:cA�|�:&�g�9���F��6�KIoy���il�EI3�$�G�N�_�y_�������l�d��!�8��*C&���Ve͑v��U`15���Vc=��o'kQ]�zL�֢����<�	3p.�&t����Q�9�S����@r��P��{���w.JΡev� ������d͜��M��|O�v��x�&�h��ͮ.���	��֬Wɿ4�~8#��Hڌhu�}Y[�BҼ� rV�����u�K�.Q�7����Y��`\��I*��b?(?wJ�~J;�~�Xٸ���j�����O�3ow/o]I�7�Ԃ���Q�&S�O'`�
.Z����]�.鋴\���ؗ���`���n-��7un�H�XP?D��-P����v�ц0�)C|]Wdaq�o��p�S���j�;�� �}O������ɸ� {�njY��o�;Q��'�F)�_�Q����B�3�NK�6��G�wϦ����L���������q�E����l�i3�j�ژC�����c����l�瑟�C#迃@�����׳���-�m	%�0��1�~5Ta�Zñ��-�<��;��L�V1y�i U���e�g�"e`�8�o0g��Kbq+jl.��Y����7���pE��;���1��*�.��I�A��%�IZE�ngc�s����Ǥ?�D�ۜ�f7���5�4��S׬-!���t|���̀ϩ�yĹ��5[?���8G���Iş��]xyh�zY�cu}D�Jz��>b�Рv�'\UB#�q��8�`���Z��9ҟ<�׈��u�����-7r+�j����yoq^��l���Y��ۙ����E��SpH�%��+|ks6��� �8��X�4���W��s>��*�����.��n�O��8�ķf���H�[!�϶��NT�d���$�_��ƈ�T�}<쥅h���3�?�5�F��S���fw�� Kg١.s>�g'�si޳�La��7}Θ��� ��y����|�_LOG�x�{�9<JMVa�{$��jⷧd�igxyM�FŎwc�
i�߮�@�ީp��u��Ǆ��Fn
('_�a�9F�������P{��@���'l�YU}L�.��a�]�M�-��K��.�����I�-j���0Q@Gv��ז\r��䞞��p�h[�_�J{;��e����=%����l��Y^9�+	������O<p�s���h6�"�{u�����1�'�ô�G����}]����A�����?>5b���n�[t�~ϊ�������
���dcu����I�e�Ϩ�,n{��U=�'�I���F�E�ȿV��%v^�� �X��օ.�~8CH���|�������ˀ� d^V}� ���כ[#փ]
,)��:ߣ��6�aH��r�_&�����a�2���4�Kc���Hz9eJ>�}4�c�"���0Y*�7���{�n�MXq�9=�-@�VZQR���h�/�{�8D��0�,�uw�P�����Ѥ�)q):�|���ð���	Gyj蓇h��4y2��b𵮐h���I�B�������"�x/ݓa�������Z�k@��Z�G��	�3��k]��0�?�6no��3��l�2�hL=Tk�A]xMf��O�|>��u�Z�%�==\����L �۳H��y�e\u����V+��ǝWBf���^Iu�_�ʃS���J�qQ&�*.�E䁶W�tp
�I_�4yx긃��C������,ѩ�N����5M��9Q������������-��
�@���l���Fr�C_���>5jRR�����XU����阬k�{�ǶR�˓�ۗ��9}�R\���#��,_wʙR�`���;Ƿ�����0u�	�Kcxbx��¹��1����Z���wv���@�[����ġ����O>�T��\�K�=��av���S.�n��%e��P��W���,��S�s�f�B�Tm���N�޾j
Yh�!jk����y$;�o@;;��N{!���
\�u��Uڢ�9o1�T/������ZZ����V�ˁYtX����h&l���@<I7\)$�xʢ�^�vW���=�3����O�a`�w���H(6�����FK8 �C��������'��=���\�OhJ�4�FEq)ԝ/��޾柭\@�gSu�̘��'n,���٤h��W���,6����;�/dFA ���#�\k�혣D��.��U��Cc�5�ARW��Y�=��O�������/������-o���A���H��QNt��^��
��<V�*��a$ �K��ۺ=�X縷��>���v�����o���$	4�pQ�sc�[��qw���ߌ��-�Kj�.���˧�̩Ӛ��B~�2/P��ʗg��!����!}�Ãl�w�j���'�K�=)囜C<���WFng�`.��˃����%��u�ձ?�_�����F���ξX���̝��G������k�K\�lK<Ǫ��r"�A���;��=�S=�.�M���c+0�n���Ka�AvS�G��m�TI����.@�C���䖦�f��k;O���k0'/*��'�K�0������;?�y�qlk�)���k�Mߧ�"��F�9��<jD34n��H�ˀ�*��Q"Z��t+�W�%��63���pѹ����H�K�VM�<C�t�o��Z�墺�
ɧ,�IZ�yET͚P�z ���O�E1/����7$�GVvT�n��F�&�L����@��j����ۢw�&)��pA������SQ1Q���j'EF�g�����o-�����EQ,V��"��vm'ME�F'���{=��w�o�~SZ���x>�+sn���3ܻPB�o,զ�/j�m�d!�t�m�j ����B"�R�<�.y�����>��V���~���̛��8ʬ�U/�AI��?i��x��o��5w�U� C��⻝C���o�qpWRNc:���v�ը>�`�XD�jh��W�V_��NH��b�1�Љd���&�&7D��+�Hݣ�� :Nc�����3&>�e [L��'���@	����K�R2�)�\���g^>U��U���Yr�|���|��ٚ1G�]C�n�D�'��F�@�� �i!�wX���i���)����r 9�F+�#T�h6X�P=��1;��uq>�9#�j�!��kud����;L8�s�&�! ����%�"�Y�B�2	��;��_�fVlu�tŷ�Ǫod�VTl6)��i,�l
Ig�6����k��@���;O�� i��V��-Z����Ih��vd� ��E ��X���-�<C���� !��n���2�߁vf��G���c[�$�3��n����Y�#�����E\{����A�ƴ�������)6��Y�%F���!P�5�K/�p9���l��IG����dc� >�����-��^��~{������r�}�N%��٣���k������w]��('f!%�;z�fCi��N�b�i�_��
�7�k��|/��W�Qn�6�W��;���&8�\�3,�%m��{�˼+D�奷���\����C74m��;���r�[,c-~���.�֓j���F ��t3��gng��-�cZ�uק@��cHjܢ���'}]����I��lV�����e�zNp*i��6�,�S�+*ixMn�!m���I��.��(���^��+��:�ax�[��wx~�_UOz��'�L��/���{@9l��X�<F�����h���/糛��;U<_ۉ���r��� ���5�V���K���3�H��ⲱ0�լ�P��m���{��!������Qjq�$�`�pM�J��/)V�p��2�wH'�����Zal�eA��)=�R1�}K%`�C����6�?�S����ߠ�~�Gb�J��t�c!����$V���n��L<�yxl��)�\���i�U��E[��ʚЪ�d���i���ހ5���N�K�c-�?:� ��KRW�pPU�)v~O@��������M�R<�Lk��t݉�F��nBLA�l��볽��]ܔ-�Np�Y������]Q�Rwᔟ���4M�3е��4a�B��u��Bny�-����/�\�byT�*����	�	�]�tC\Ѩ��a&��;�͸x	��%���w5�������5��W�8p.v���U��[/]旷�N�)������R�u�����t�ұ,o���KX�ͨ�S(�\"��c�n�㯩���ԡXr�tS����eޗ�Β�J��C`_-���%�}f�iRM烤��.{(�J5��	�d#�
�@�ݤʭ��N��Z�A�X	"��cMb�H��dcĽIdt���c���x��Й�|�L�n� �2���WJ�6�~m�#m��p;{c�ǧ��]�{I��y,)�=<� ��-22�i�(��ä=��ܰY����om��@q��ޞ�T]t+#K��v�[��]~�Ud���`�k.�����T�x]��hS��:{9�nA�K+�R>	�eEl�Nu��V�<R�0|"K��q��U?�\�Q5���zb��,��0a�ݭ��5z�#
!I6�����;��{L�k�a�Q25{��e�wH,R�H�D�h�[|	���=%L��jm�����A�'��ҕN}��"�V��a�>2 ��Ҫ��CB��z=�� j���ya�&kR�/ooKm�t0� @�7zDl��l��B�wHF�\L��O��l�Ko1�P�~}HN��}�"�.(Y��W�x5D`���EU��%o�F��f޴  ���y9�#7˫��d�:��g��t��(iZ�`fH^�X�������]K7=Y\��IE]�[��@�Q�@��ŝ&RYJ�6�\�I��X�/jjN�$W��ݺ�/¯17���d;x��D��@���9�t�����A����moF�7�7��b+I�߾^�Z��	hw�=�M�o�B���`�?��茶���h�rH�\p�[�o����ܼU���|�xQIͶ��_EM4t3�7��C3Dr�v�s�����<��n���I��� E�sU�\���3�@x�#�[�b=�-@�2W��-M@@����������})��^����d�ffeZ<��5[g��A�/חlO��<��_<�g�t�̹8�������䊨��\���H#{0)O��
��\lݖn���s�!�\�A���7��)�vj�C��^��\��Ms�f�lr����,��:�H�7a�o{��F �Q#ܟe�aͯ�"��]�?�|�z�>H��=�F�«��O���jR)��GH�����{D�/��Y��J�(���B	��"����^�&|u�Ҫ�	�] ��bi�q;*��|Q���|$�PD[G�E�Ւ��*�z�����͸06�E���q����l�uƎb-Vj��i̬��XX��V<17[�L��mh���9N���uj��5g�Q�J���q���@z�k�
65n4K6M�eҍ%���	G��E�򾫠:`����R9$�'�~u���_�>�>u��ܲ!9�ȩ6ьr�>�&��ۗw������[��\J�ŋ;�w4X�{��}��Y�U6'�L��CP5�#�=�3��$�0�>�O��/�ْN/�=�/I6�9��*��թ0"�kjsY��+��KY�C�AB�❴�73��wܳ���3b~�Q-H��
s<��C�����`�j�u��ؠ��V�^���
�$3�>0�l�/���y���&;��J�֨$CS˪;�� ��]~�d�2��	F0-�Ju����qjrF*�N���qu�]˔Y��)����b��
.��i�r�0���������&��9i_	�Ƀ�J$;9�w ���:�8�Ϝ�үo�u%
4���� @�.�_��+���-[ �6�P�9�,w�I$�C�ԉ�n�)`�"P��r?U�����%����Z��\�ڑ��Q7����<���q��n�hn�}��sF	��mئ��r��] r�xm����NF/�Z���,�ԗV�z�.�K��D_�^����}�T�=�4��er� ������ B�83��B���L�"�0����v�jW1c:�����II�������x�M���FQ��W�����ȱaK��'OE�l8햿N��v�&ŋ���{X�g �����^֨F��F>;����?���}�hK�����آ�yh,��#P�O�����"x��_�[-����(Z���F�t�x�c���He
E�͕�b8��u�ɭ�����*�YW�o�S�y.����N�ʸ9&�ˑP,�H�N�y�>Q��+�����}c��W D�|z��h��!jӨ�����	�-f]�B�X����V�l��]q3���U���^�޺�ٚ�km�f��l��Q'K����=�����Ugꍽqo���$I�e�W�\U�ݐmc�����7�<� ג�2�!x-���_6ate�$uHj�]?ۧ�í�A�A�Z�*��T ���:2@��N�B���,a*
�����a�U��]w�ԯ�iS[�p	���N�:��x)�Ukw��U!`�
��椭�7I87������<��p&!(ե�G���|#M�Э\A����G������z��/i�	��|& �
��/����p"к��^�'į�,Z^�kv�Q��y^uT�����WV�S;���3|w���
֨T��o�Qq�0���`8�_�0hW�����;w�u8f��R��־�����\�ͻ�B�r�e�1�qjer��� q�<�?���x��/>R�[xK��BZ��u,QYb�,Y+��o�0�T^	!d;ٓe��P^�}�i��$�c�0��jy��<���s�s���=�޹���d2uD�y��P�[fVU �/a�rh5#�L4�zE��#0�V�p��L�az���К��!_h���U"������3|��#���
��<��s�_��:��2�n��rʳK��3�Z�C�Ip���Ӓ!rZ�ּ�st��UՄ�w�ӝH�P�;&7���[����%�U�s�~<p�Y�aq
O
]���-��	�<�_�[��m��ßj�V
Q?��q��3>���,9�iL�I��~˸��b����^�Ѵ�����n��/wiZ�{�+<��Xf���j]:�x)�����p��|�Q�q��(��a���:r��i���#vh-0���Ǡ<�:V,�ʀ�#0_7&�����*�q�]�F��r�h�&�����T�����]�u�1�<���2��7�>�{�Ԣ�c&���	w��4�J����G
u&.��M��G����ڎ�6�صZ�EN5�Ϭ�%����)���տ׻��䶴$~�l�޾��m�ꋰ�-�Q*g�<�LX��>�<��m�y��޸���e��]k~~��28��@�m�X%gZ��lp2�x�^s�G��(�ҹ��@�`^
?�?l'�#t7�o��;
~s,c��F�ZWՎ�����3��fX�D�0���������2�fB"���|�5�M���F�����;�0���5u����jaч�����@�4�[r}��a��q��Uy.�R�vˤ�F��N�Bo1wϡ��3}ˌ��}}�ã�;����hR�HE�%��ʔEig&���0�[QͿ�;�W���؉WW�S篇���[yQ�a���}�t[�sY4n�NUU�������L�_/�o�Z�m�.�p�����Ғ�ө�1�,��"���%=w�������t�e�m��V�_�܁gV�)Y�nח���������q$<g'!Ɖ��l(�>U��i��Dm�ٲg*5i6��XLM���E~"�_�E�e��TMl���s5��I<�B�w+��c���<u����V�3�:���Ū������
o{ԕR,��q��-���3��}��8�ޮ�yʪ}��nHt�\�.������#�^�W%��-�n=9 8,&�M����YP���q{`>.�g�8�S��w�ߙ�q��2��򓿰Ar�:���fN�"a�L�Ӄ=#ˋ��D	�c
� "��A?-w���}!#�&#�m)�r�j�[\�)Ύ`�!�2���h;��;M"��-�K��}Y( �H�&���7Bύ��S�V�<'*Y�M�sJ0��F��~G/����^|ǧ���3�FE��ִG��V;k�3�i������C��+#�O�g��y�-��$��
�R������4��v�Nj�{@_ψ�uR��Q)J���>߇���r���K��k��b"Y��Wޟ]�, �j�^�F
�姖�z����殸ڄ���M.��j�`{LC�@L�N�D9>��M�j�M{pK6a'��m7�9�!���E�g5�*��.ÿ́dW����Ry�P��S����_����K�'0������}���<R�"�R�ղ�\�~(�@�c�ϐ�[�Z�Y0��X��`&nmWt�7�)Dy��Qz�0R�q=����:���EL�Q�С�Ɏ
�ӕ�j�*��{��y�ܼ\�e)ߴ���W�U���j5���3������`��\]'G_�G(S��BN�����_�PQl�,;��)���Nr��n�6����:mf�}�Q"+`ݪ����M)���(�nӃ��A9D�Y�%[Mx���鉿 �o4�z��x�1}ϕ���d�:K������v}󋚛�%�%��i�b��;��rЉ=xp���½S �����$�W�0��K�)�(��q�������{�47�V��_��UYc�^��Q��}���G\���e1�c��0�&fͤ�X�s��ۀ�j3��-7�"�(:U���S��U�8~�O}�_������2�mKd�<�D��T�mu�*������ot� _كoA��'��A�ӢsE��!�S���u��[}�X��¥Ԛcjuew0��3�ja���E/����C��c����s�~���{�;�%���k�!�^��<���!Sno��)x�e�,B[���ja���۲Նɪk*n���T�X����1lenͻ%�`&��.�
�VͩpEXv�͘5��/7�}�l�%�;{�q���!e�ir��#��3�i#>�#��(Sޛ҇��W�+�X2��"j��B�,�%AH+LUp�����;��(�������"TmY,��KC+^V;uul��Ի�n���w����Շ�����r_���C��\诫Sn�}��Z��Ǎ$7�?��y��g��!�{����vg�w�󋲎`H�@��t���c.s��������:�ё���K��*i�Mۙ{+h)��]��Ԫt��T��%��Z��6'�>�6�����;WQ��:/�*�~��+Bg@�i�kԊ�{�ڤvt^,쭃������ٽO/0�04˱/9���%H���
ѷ���jҧ=���$ݩ"q)��0����=q�#�(q��f�(��0B� 2/9��Z�@TYp,z~+�E�/8ܐC�(s���NE��:��ͬ:�`�N@4�v�p]��
Ԅ�%8��m���'�G�<�j����یa��#���h��W�� �z�x��3�S㽾��w�1!A�j����$��:���K�=�D����¹���3��,񉃕N:N�}��O
�d0�;.��Ka�B�C�"[R�o��B-J��'��o@�r,��o��s�7�Ô-Q�jt��/���c3�1��s#�j�{������ ��:�`Jl�r�A6�N1s}^W�o�*��䉣/�p)��@ruڃ��<T�?t��:��w�SO{�y��l��,�ʥ�j�L�}.J��k��/�������ڔ��b=8�{�� P��z�����c�X5������ݾx@��g)��KwԿ��ӷ'�"���θ
m������G������[�|��&�5Շ�c�<o�1������d�3�׼���;��ŉR/�_+i�y�3Q��V��솒�~������`0��UmZ^S�T-#f��9e�3zG�� [�A�ڷ�G���V���*lʆ�z&L�냶�v��t��ݫ�:�6>���6�D�:��d�xF4�C6>:v�"�1Z��j���@X|-�� %�~�7��H��&f��x���Z�K���(�]F]:�򌢺��w^�Z�;��%ݪXN��٪mT��-ۣ�h��.��
�r��1��:��I�Y�c�e5���v���$kb�}y�q�Ɖ1�v�L��r��p�|�s,on������0'uo"m���@���< O1��b}�(��b��Rg�Z鸡����S
���6B��q�Mȓ�<!O8A �DqJ�kyYW5v�3���ؚ��NQV��2;�(����>�ټ9�.yX0�]��cH�s?%NT��Ek�Q��`VH�چ,2No�/X6���j��>�,z�t�z}��.n��n�^�=����PJ������[��t���IP�@b�RA�R�r�6�ڍ>��{���>�����83NO����ʅ�7@T
�4*9[z_��Ul�Rɵ"�0e�{J�[󒜳fG�<��VZ�|ɱL����C��|�g�I�x�0�plt�>����}�K�Rp�"G�Ksw��3m���~~=9\vj^7����8\�z���	��5���=�CY��롵�G�<4�=G�.7bl�I(5��4��zK�.a���LD�\��K�F��_/�,��tuE�%�)4��Yĩ�����ߢߓ�!1	�ۿ׹�x����*����k�E����`h�Vq���OF3��u�]�Qec��>Q�����Y��߷U���3��#������C��R��im����u�s�YV?>0��p�>�,�
UVWap��=lk�Ya�^�������˨0��@x��¸�bd���35V)�Kv�Yg�یT[[�����}����᫘�4�l���[���8QKM+\�0y��fЮ.Kk��E�u����߆q����=��%tY���R�2W_�sw(p�ڸS.k���M�-q1
q��!g�]��ƫ�))%����nC/�[X>�������f��Ɯ�+ه����v�/ɔ���1�ٜE�Wo@2g@�y!>�F�J��9�ܒ�(�`��ݦ���������d��ۉ
��U�q<�p#v�}�Ǿl���{C+�n^�使g��!��aE�t��-YlbKπ��J��lz"GڦF��z{�&|@�W"���C/2p��a���(��#Mk�ōX��,�z�.�TT��3��X���Ԉ�}+4V�3�56A=��5���Z����QÙ���ܷf�IM5��c�f�6���T�k��!���zG�zb��xU+�{�=�✻D5ŉ�K�6��Ά�3�>7��K��m�-�T'���.��H\Gj��Ϗ^oØ��7&jj0�����D���4?��4��X����'x�ݲKr����5�bRZ����gX'�m32hӤ��e=�a�y3#�`��N�v2Þ_@�������H�%���x�2�s9~���:U�AF�x^����G�1����(<���&�O5ٌ����=2Pm
Mp��8`�����ec䀻ǟ2���)v�d���:�ׇ4h�1��X {���kI�����ɯz�t��
����<�%�����qf}�=�G���b����v��U!��g�9����Rcvd��R����V�]W�a���t�ap��xW���^ޖ���Rۉ��K�ځ�21x���&�~mcc��W.�bì{'�3��aϰ�飋�8<�/d�1��5��Z�V�`��$jg	Y0ה6�s����*ɟ�y�,��31��b��$��m����ǟ�bE�j��q-��Why۪�̖�e R�-a���2jPmɾ�z(�O���xp v�I��7�Ῑ��[�;g��Mm��Nr�<��Z�Hus_�H��uW�t��Q�(i�u�;	�ܽ,�b}8Y�D�k�Xmk	X�8+�X�b�*���*��GgM�"��Ŀ�@"-�u��L���GrckuI���侏�{IF�+Ǵ�5�1Qc��!�Б�	(O��� ���1Ο{�)�X�;�9�J"����w�zx���-r�n��?@��w��3~O�e��2�IE"�����+���t��zq��8�����X���~�����K�&��ʮ�C��<Gu9��}v��?���8Y�K�G����+���F5�}E6�'�R�qݪ����dЃ�W%�*Z�������Sg������|���?�X���c]Ϩ(m�m��˴��%]XFG�Ȳ/�r����������S
�XN#�����K�[�����I^Ώ�>�ȼ	�X���3T�N�����J�7�u�چ�u�"�l~������К �ǥ.�1G�o�u��=H��n`g^V��Ӑ���"na��Q���Ylٷo�Tį���VNz�i�۪U-���v/�_��fs�b��ɽ�h����ó����Jq��~��ki�;�l��7n8���ߗG�}f�}&}.��?�֨�9���6��	xB�I5��GlQ��+9^.O��j����5m$w.x��v�c��o��NЄ��r2�ﰪYF_~���^�X����A�������$�S��N��Z���o��}y� }��8���b��m��'*�q�Q�\"���)�vc��� ��ӑ'�'�p+��D���I+'�K2,�x�͘�!��	��|�\tM%���D�g6[J�V�ĎGl�����+Y|�ӓ�s9D� ���g�"���E��~��1tm�$��g�dw�m�ƪNtzEԧE����+��_�b0&��ei9�!��-v�)�D]z���X3�r��E�w`6�c��5�4!_�T���.����w�Y�����7���%�I��v�B-�÷?;�R_���	���ON8�1 (�B3l�������;�Z��F��2"w^3��ud�.�"��i�k��ꫪ�~��wY��!�y��������ޜ��M�9���R~��?�I7-�n�y�w��H˓g��[1	�?7��3��3��Q)������
��3��� �/���1���c��%4<F^�}��9��C����_!HS\��������;n�-m��hi�z�Afkğ(��R<��C��ɚY�ߓE��!����� ��R�����\�f�N�M��g�\!�8�O�q����ܫ��S�nL	i!���Y��P����٠��z��Lon��������)��1���1�c�H���|��o��H�v�Ԍ�~�)�\9��<�$�!�,��96n%8�������e� �Rz�Q#��.��l�kt�E\N�������?���Cey�{O@q��Ε&�����<q�����-����a��q��=�����LU {�ko��v����{�=9�ۗ��?�YRd�N-K�T����B:)x���p��o���E��"�%	fϟ���-�t���G�Q���Ѐ*�������S����*n��F���=��c�\��~��f�+��Ζ�Yl���>J����*8�:&8�6��ot������Y������o��V(pRA��m%��W�`HN��J2��@�KU='y��i��9��;I/�~y��w��z���XF��k�u5���_�K�����W_=��{G;>� v�@����9]�cC7q��`��0���x��Q��&*ܪ������jJ��{�[����*���8/�Bf��=���-��`�\I,��Y�I|�A����M�c����V�3�Ԁ���2V���jR���Ԑ����J	��G���)y 0:�߃��:�}#�=پ������qb��]�a�t��qC�\L����uK����iX��8��z��/�[`���YeҺ����Ƭ��%��Z�M��H佧�t[���[�#��v���y���%�Ij�r��u�/M���8������������p���l��[q�~�v�{@O}\'����ճ1.��o��^q9gPE�W� 7QO֤0�Q<ǬN������L� �\!>��٤Dѥ�F����5�
�_�rv��/�uk�p���J��=�{ �annȝ�<�ȳ���?~�Pq�s�4��U�Y_��ߔ���ڠ�t�[_Y=�?������	���4��`�oF�>Q�Ŋ�I��Q��Ʒ=�o�{Ή˱�����+r���滩"���%�?:O�O���G M������7-ң�x.I�/7���\�J3M*=�dN��u1��s\ j),��Z.���N��SJ�s�z�ۭ�4#jc�U�Q9����a�|dh��+<��w`�2���S�;�6��՗~Η;O�s�}#��v�ɑu��Y��āB�o�j�&�"-������9�P��`L���r���#)N�p?���W<�{�ͲD�*9�醁��6P�V�IY��vڶ*��ǡA�3 zv�7&vT�H�S�%�.jvO�{�y��P:ac��9/�e�M���p����#��g����ob� bȂ�[�٬#��S�;O�k�BkQh��*��s[ �I��.ɓ	(���*)�A�H7'Z�_� �k����0�a��p�ף�4ˊ����@$�*���7����� `i_���ɕo��4�1��4X̓���rjH��>��9K��s�`'����f~�� ��$���G����tN���w�a'/"Ia8��S����V�!�iO��n���:�,wk*.��el�	�� �7JHhի�ʬ������e#Cb�)~�3e^`����O��ä���%qI�)��[%���R� <��~@\���u�&��`f+ň65e+�D��-͊9���e[�5���b�Uc@^��4Ǽ׈�jc�Mv��;H�����͵�J��х�^3�V����Ϩ� �K㮕{����mt�0/{/�0~Q����JvY����}u��J��� �Z�p���«�ƻ
\�jM��u�@����������H)�pK��Y��l��~X��{���٩��n������@qEBe��2_#�Q贄��/����"`;	1��nޜ��[� ��[Xi���v���ѧ �C`�����������2A���e�*����і��ٶ�Py\1�
'H�ֶ�6���� X����P��qc�->]�Ȫ��T�Ũ���r ��<.(|�M��|�s���w7��fO���=���#�	v���~�!O�qZ3!M� 2�hR�����c�E	�V���%���$�TL���h�̤u��	"�
$&c�;�$�~R��d��)v⡢{�;�Z�@����������:K2����EE��W�P�B��b������=0�km�����S�.^P��fr)}�R�&H�ʤ�����~D.��q%J�^�5���^��щE���K6ɞpqȘy�T,�-������/��T�'O�_���xs����-����\��b.�5iƙ��b\\*
�m�h������v�d}+��vZ�e�#d��䢻��
�){��L��:�-b�l��߿����Lb�D�!z�l�R~"���{�������<��{�/Y�ɶ�hR��P�{w��A�H�Cr�n)`�RW�{�eRUYS~9q���aK�O�S@��1��.�ր��Y
�hz��9�;�C���#�F�� ^3|3d��!U��pY(_�;|��sqN�\������
t�)���F��]�_��I�X��4|����Ů���Cy�.�~%h�O�Y����7:�����k5}�(�.$��� ��8�iQQyAo���`)�M~����r�(s���{Cˬ�|P%�~_(U��*k�.�9�[<�<?���7�a��;1��b/z���?
Z�Ī��{�  �k����k�ju'����ٻ!�"�5S:;	R��[�-b����������_	'��S1���.\��%�;>�`c�+�`fg-PX�����G9{0P�E����͖�Ǝ���+$�>�_����G�pe-л���g�	��{�(9���tE�UbF�
Y�?tP�jo��C���E*oG�^��1C<)�@��0�� �W2%�����dj ������E�"=2�@WA�B� �7���.��GA�wTO|�:���Y�F�5b�3��#7�A�� �Kl�66�C���\�4Qt,�����ц��#��.0x=�u�4H�/-W��^�R�5ۢ��~�z��������&qw�s�(����?�s,�we>�=ê>֤n��P�C_��Zv��u�Y��۟���v�oVt��V�};}�Պ�	����I�=�<=��.&�`,x-��m�}Ԉ_�.��}�L~Q�2�(j�tD�+\����.���52N~��?Pm���׃�d��X���Wo[EAޮ%J*r�Ow&��sV<����f���a��PWR@,"T��vtŢ��z���G?�dU�q`ͅ��U���ҵ�I'G>�JȼF�N�n����d�W&����n�xD�K�C�O��qw?)*�BI^�ɍ]
�?�g�-@�`9�v�ۍ������:Kwn���W�A<9f�1w����>g��x��H�8{;U�}X�@���E�/>���o����V�k���DU�Ug"�%K�+�}]ED���U�~W���B�j-g�Ɒ��*B�t���3�"F��8���D����կ�|? u>��R[�֐��?iq��`*Ef�V��74�-����w�C��m�\�Ĝ(@�|�W�!;��="��p�G(�*��6��]�	�����~����W,��U��P�i�Y���|���������A�6�au"�DI<��\�3t1?�����}P�,���� l�2S�F\+�`��; \��ۀ��T�EѼ����ΩL}���I�z�7(<������D���r$FP��v�&yn+$�'�D�C����f����ީ&7����b�!7)tX�^�⪘�[�(��R��9_�\6ʩ6�%\��ץ�|�i�ƈc�$ζ(TL��Y?�O�s��;���XMkD�s4m�B{B���Kޞ�v�*�Юj���S�k����f1��Wu6wbx����;6�M�G"�T��6������l~	�=�t���D��6VӴ���Tά�_N�% �ݾVRb���N+r�t�I��u�da�wvy��|x}0.w�����=z[�!���a!{��? ����BeB�	���!�B�ƫ�Z�V#��j� ?�|�� �P��$Ue=��ό©ފ���N�<6'��qϯ:��,Yʒ��b���` �<i��
����p�D}���/E�� ^�f@�?�}A-��c�����z�9l���R�f�`Vc;9�E�G�k]��p���R�J��`@��.�쬑Ju��ȁm�9.�9I=z*Q�f5�W�z�5M�I.u�ZE ���M�Q;�.�k_����kQ���U�l1�H8;�;��#�)����#�@{���f���� �9Xz���.����֘��>��3�����e�K곁�1�s�8o�sY���7�r�E+�$��_��ӯ��ѧ������z3� ����ٲ��P//��R�����<u���H����7���e�v��|B�
�޲e|t�A��y��4�K��3�$��7(��;��n{ '4�_*�x8Pùo.�V�p�w7i@D��"t���,�BW�5g���.�w|����J�׍7D���R.`g7<`��]7�rF�B�ׁ�J�-��EV�U;��h-#u\����p/þ%��ZpH���y q)��e���qk}y�GO� �u]L��߱_\ء��Yd�<n�i����
lO�2&�b�)���A4������f��W��� �w�X!��4��rY��@n�1!�AW޶E�cE\�S\��e���A�N���Sk?�J*:�]��4��%vn��z�ŷ5W� �\�z�
sݗvC����t�L|�@ L�k��L��.��o��s)j�l�%:�46��zp+d嵼�Ţ�K(o�H�L�V�z&���[�Tǉ9
xѨ*���]�ʷhji�g��"����.@u�NYR��^lK��x�xlG�vVz1.no�cI�hE��v��\dYeY;������$���y��g�(�j���tU49g���*fg����q��gQ��C�s5�����}|ڴ�]�B��l�����x��ܕ�T��CeOY;`�̊��`����Hz�շ���\��ό�Ծ�� �!�.�H����?\<O�lM3bw�d]�<����Evw��74F$pj�w`� �M;��!l#��;E�k�U��>۾��R.������J�~���X�Z�U~~Z'��BwxN�iÝJ��l����V�)�ۯ�'2��'�q���\�{:��ZQ5[����s�M�^2$�k3]W���ɋ9���𼒵Ν�9Z�''�	*��K.�#ͻk8��,��t8���D���F�m�z���ƽ89މf�u	)�}/,*7 Ҭ.�6�:g}��w��S�ή{�А�x,���f����*�B��/�w���ZZR�v>�3�:*#T�u��;xK1�"�k��M�H�wZ�i����0�⤃FoP��p#3�
��|�L���:�l��%[�Ky%�냘��e��O�i귇�O�Dht�P�/~�3l��B.��RU.��~�řk�z��f֔Tu� w����<{����>��1z�g:ŋ�x[R�<4C����b`(8s:�H�;�@������ypG��5��X�6���k�1�|��k������m35�1|�e��˯Ky�ݍ6�`w��{td6o�'�}�fB�^R��Q,~�k��6�H)��l��?����v�A��*��g�s�b78���f��Љ*�m�Vժ'�����SZ��^S��WD�ƛ+WT�`��A@ ���6��u��w�M~л��a_�jpB�Y�� �ݏe��Z�0E^��7�@#کU�ϣ��ҿ_��*����_$'һ�r��}�~��M^P�C
^���P���"���J��\�^�૓e�+��B�f!�u�ޗ�eUt�M�7N�&�@�.�s�v�уD�{�[��ocB��#Î������c�2�q�ȃJ+d|]�����9�+wb����c��� ���M������Գ���sg�Qr,~}Sе/�g�+P�w�f�8���-�V��W\���~��J������n1�;2��\Y���T�+�t=�u5{iuX�����$s�%'��e2�q����۷*%��������}[2��M�Y�ڛ-�֓���0�w'�hR���,<��1ԋ ]2G7�<������F�������}֩w'	�����z���;i�qR.+���e~q�в͸c#�f@��Z�eq��f۱�+�������B
|ܠ�{�c�U��.\j�c���Ä��\��k6nQt�k#�ً?Fn�~��o���̘��^q�}��� �'��p�^�W+���4 ���h��͝!و
XNV(Z��蓟��~{'�'��ҷ,�v�"D�+Oغ��]��-t�D_R~�q�����Ph��N^r�_��-e�J�Uڢ��r�V�f����'�z#���7�@g_5��� XhKyHQϣB�9�Q~����i^�c�b=�J<>�p3�y��>����~ex�Eb|�+�_>���p����%@��?����~Qww9��\���3�� ��Vire틑���$ε�� ��3<��Ι�k��00�}�Y�]����[��4-\�
[��j���X��
1Vo�	�_�*�9F@���4�I��p���i�x���*5��g��Y�k��蝁o���5B�j�{�`�F����j���MjGE'WH�6+:��CO�F���`�&׊v�GU��@�������@��tiJ}�~o��IoIB^��Mp��f+�C>�3��ͨ!���J�h�m���K�cǑz����3��4s�����lE�Hu�f�md <�\A'�L��D����{w^M���g��-�P�֗	�ׁͣ��Ђ��ǂ���.5!~*Ë�'պ����q}�
 �7u�`E�M^�#:�n*��G��2�m��~R`5?ЫX�(�5��X�<����c�E�.���t1�&��,�d�`���k3��6�*����P��W=?�ƍ� KrZ�ؿ�����ؒ��I�r�q��»D���J�tM�b�<�j�mp0�~>�vXΫK��8aH�m�z$UN��~�{&um�2��Cr���1O��6pj����X"��o�ޯ,~R�;e� �l� ұ+���t�⢸�Y�EE��0es�qYVHw���L�n�KT*u���pԠ�:�&@�7&u!t���$��\[��Awm��_ܺ'�Py@ɸ����� �1��f���e]��_�(kR���n���FM����y`�~͛��}����|�F���޵��2��k�,�@>I�"��B�ǂk�#F�*)�bT�A{	��M�%�t���4�(��mG�-/��Jٗ}����D�wa���W�`�Uxb* �������*8w2ݟM�{����l^����$f�933����E�z��O�I��
j� ���5[6����+'���$�x�r�����qtzkmc�?�DuCf�&F^�sO�rk�s'O����oG�i_$��|��W��v=��遅�S3�FZ�9�d1!����0�U^(�"�UA�H>eS�H���<�tQL�|$KeZ#�T��e}M��J������i�I�x�C�cQ������P��!O��J2;�VSF�ٱ��ݜ��"q�[����� ��7~���4�نϷ}�O]���)
a�q�f�{6�Q<���y�����g��S�FnI����$4�	B�[nA���Ěl?�&�2S/J$�8�]�v��v��V���p �\T1���ў�4*:�vu2����0 F� ��Tp,��[S��`6o����buG�ؔ���$(Q�+l�*���M��Tu̶�G���'���k��*�0i�`%�F��#�D�x�0�gia�噐�֗+[�1��ئ���+�4�r�%ǥ*��	���_ȫ7&�5P��J��A1*~���I3e5�D�g�����lUߊ��dWζ����$������+��7��/m����r�e�����sy�m��]/�70�69e��t�O�9c��B�R�����jچ��mZ�P�/�o���Km+O�4Z���|*&c5�w�Z(��Uږ���<~�r��fN�p���`0����U�{��v�i���c������>���_!OZ{�(
I�Z]cQ���5���-v�:�����g�W���
�a�U�{�Nw�{^��e��aMsJ�s����ӊu���c�~\s�yJ�g���&����K�2�&�zEH5):RǷH��K^�>�P�����~B}\���D� �� �����7�N��}_�oo}��$��V�+JJ���z7i;��I��j��-"x~�|-���HgbnvT-ǲ��(dK{�F��o?{)@QL��\�]�]9H��'mz�+sk8�j�%qE��Ee`���K�RڔF�5g��(mu퇹F��i�-���v�o�yq��-AF�r�3s�E��9ɪek��g�SY�,s[#�*�����l4ٺ_�$N�4�c)K��f�CF�/��"��
�6�4�W��+��(<:����u�&��I]�Ď��0k�}$=���/����C-�4�7��k�P���`8��8"E���)�@�qY/c��>�{A,?���f���4"dǼ�o�������l��G�������?`F��^�Zyum�O4ױf�'�,����~�wCUG�n�Z�K��K�~��+�YhQx���D�8#|Z����cLK�����o�K����j�]6Z�F�S�G��V�c֝Ȥ�WQ�'24Q��rKԷ$Mθ���╗�C�jS؋âق����v���cv�~+�0�}v�gE;��t9g=��is����<�)����2`�fy\����|nU<��_H��	:�\H Z(Y�$a}�!�c�0�Q-E����W�$�:��`AE�+q
�|���:*�{sb��Zxf�Rr��/\d�
���7E)��1�@���.T�Wa#3qp��&8�������E�&�%P�b}i�5����rη�N�	����h��3��>j�^�\��wB܅�S=���W$n=��1;�r�w�v���M=��e�:���Ҳ}u�Tq�_�F�_Sj��dٽ�Y �?J�'��=�1D�}��{f�z��"�������k�f��s�ר魵1�j�j�� ��P59��m�D:�3�@���q8N�w�� WA�?@��	�'0=~���މ�|ڭ)���
��v=�@Y̖����Nn�ƱꐑZ?#P\��	�jj@�'*�ݑ6�غnW���Z-D��	$�������]��݋�Cr#�T�{؃�߮�yX�y/�a~���A����)ٸ��3#����-�a'԰,�)���1�K�n��r��4Ɋ�N��@�'n���b�E�aU�������5�"&R3�H�z�yᩎ�V�soO��<��8��>W���$�q�pn�룔�����"&0J%�˱Y�����>�Qq�r�.3������nD��`��$+M�7#���"3�B�xV���HbǞU������|��_�yա>�c�@h�����_Y}�ݻ�A�]_���H���Uh*`wN��:z���롃<��}\�f|���ve������C�7&����_����EU��xCС�J�Lm���+���`�/�
��2����k6[��;�v��.���{�#��֪�h��K�Jճ�[l��u���[�2/|�9�^��/��9]�W�+@變 &&���o�ĖU�h�Cј�5����l���1j��W��A*o�'�w��T���")&]O ��bm����[_H"����b����lq�ܕ�J��@�Ow3p/l`�!'��aW�����XX����x'h������?�Y$�X��ɫ����v��%�y�z�Ԕ���D�a�e=��4wW���O�e<�]/�h�|���2ooƿiZ:>�m���pN�+c��-/V�	6
^���͵l#jA ���$�z�8")�+�i�r1Z-����
�cB�&a�6��fu�߼<ԴUO����]�KO�4';�&�,��\r��'J!*_����Ư>�ne���MV!�D�*�XH2�vo�V����a������M-G��:��.>�lH��z��o�[�X��=���c��ܧ��M��]P9_p5?m9&<�(�jv�J�҈P<���㳝oqk[/�nLte���|�k���i��f�jI��6�X�Ja�gw������͐ �ӏ+A��U��<V�Pg�XLupO~'Dc9\�k{X�2m����(Oyq�,��6�7Dbk��험 �b��~�$v�Q�)�S��+��PA$�	��Y ����&�Α�oOl��7d�_̩�f�;�I���G;n�}G�ˏk#���W��A¸���:�A�c,�`�����;! ��F��G�}}��h���A��î�Q�\�B�i���Ogf����vn���렟�t�����M��e}���F�k�}�8����ҝ�]�iAZ�{t#���������������b��8��y}o�v��wg�tj%�{�_���O��3._i�L�[���Q&��[Gz�be�MX�/3y�P�s��e����;%��7�@��fIs�,���>_h)�:ʃcĐS����>�Y��l��c��nlJ��D��� ��UYIw�̂�����L�C$�v- �ȳ��"�2e#3��4%�IwQq�� 3yX��Z��D�$g����p��.������n1o�z]ht����n����/�7&cN����Y��%q��2��9���r׶B�	e�9@��E8�(O�+��0���K����m��#�m�����l������S�X�z���q/�
�:�4�j���H|����I�Ϲǖ��̭7��E�hTr,�PZ�I�@�͆�2�q�G`��߮�[f�������:�f)(?�������P��t4]d��p0Xv�ѣ�Y�Ө]�9of,i�٣1��ʾF�/0t�^J��w+�m�1�ʬ���,����Ԫ�Ȳ��=ʕu}.�ؼ��>ڐ�t`�"%����X��X�Y+����$2,�2�`O�thN���-Y�,o-���_�	8����l3]���*��CQ�%L��H::����ͥ}Y�Շ����	|'�����kq��C�pW��s�����eJ���o�@0"	�g�cɫ����._L҃3���}��,,,�����v���R�g�\���=�zL��5ɲIΥ���gW˒�VR<S�g�Օ{��o�s.�b��<M)F���e$̭�c�hЫC	��u1�<N�0�G��!�M����N>�i8i0[ϨG��j),^9)L֙����^`���Ե
'ݏ�F�C9��mKf�i����B�/�[�;f��_�hC3c2�.��tC��ǝ�4�3������0�\[�ˍ�/O}��e�����;�.��Z^�v�u����4��G�AY��n�7-l��=c�n�T�Dc6�w�Xߋ�~���@���m��@��$r�|��>*�Q�2u��ҳ���(�9�#�?��-g�I�z�C�2b�C�~91��-��k��n]{�x������{9lT�Ջ�ϐ���r���Hð6QS��g'�����ٺ�>��U/�$�;�J�!�ɘ��}󄞫�{9��w���p�<7��-���a��!��R���Jd��I�a����<e� �AK��!�R�y��k��e��#�Ͼ��sT��u�p�	�=�iz�:�#�s̸k��&)R9�^}c�J������;XyX��;��Wa�#͸U�V�u+z��G����| �3�j$_B��Ջ�@�:,v��X��Q/��@��Eފ��L��)Ί^��RF3�U�����Og����lg�'R��j�A�mj*×y��S�d���@�:�^=�'�ٷ1V�⒕a���E�����ҍ��;.[���������7'խ]��;N�ۚ�<*F�p~�}YHd���u�@:--g��;���������扆�i��Z)��#;��{?����>�%��4����<L ?�di�ޭ�	؁ڌԧ	�����U�Q�^}~6�'���{ڜ��	|����y�d��A�f�6+�\O&n���ܾ�:��p�}[=ֽy��b-�&9�Q�0ǅ�>+^g�6��\�yy	S�XB�����nN~S/*���D���O����ox���q� ��^�*��Oٽ=Is�M�>��4����.]x��]��YRY��I*=M��G������z�\�e&K?u���
�/^[W�n����b�k}군�*���R�c���NI��&o����C�וY��к8���a�� ^ן�C�$��c��`ħ��$�ٚ����.1L�v ��c��^���:�����lh��m����̛�^��Jǅ8) *��ᒅ����^�|�]�{!�v;·��Ƙ�?��g�����%'h���v�A��� ��	}9L�hu�@#�ƿ٤���>��f�\����w6�n�F_!���	�Sܸ'��<TǮ���Dߣ�׉�rp�қ����^���ޡڴӌ�#>����u�I�D��~������S֎����N6����jl !يB��e�-��{��럃v�I�C$*�����
�m}T��Q�ә~����MEsɔ�;zn������٤Aw�âe�ңu�1r�C'������}�XƇ~�yvGx'��w~�%�Ҵ��8�V�;�|��CGq�c�x��2���/��`�׋��{i�p9��Źn��W�t����N,�k�#�}�R�=i�o�R��p�7��̖��k����m�-��5q��ҭO ��;���{s�ýF|(���洭N-�����l�_���!��
���e�W����N�`�v��X6���G24�6]3�R%UP�
�3�O|k�*4wWP�H��C��4`7��$����OX71	���z��.I����uw媵��W�	�����"L5sn���H:>HNZ;��.Y[��:s��NJw����v��f"����߯ŵ��������׫�>���� 4�~[��;Deo���>�Ʒ$tAHȢ�E�[���W]r�� ݀.���Js9mfˬ#��
)f��HoD�57Hgz�� ���o��D��g��z�*�H ������6|	�x��
=�U�K���olQNq��Yϥe���b����̄���7����Q�'-IE�f��_���Q�Ѽ����ϛ���Q��ዞ�wS�~�{���Պ�u=�=R�<�چ��og�B�@_g�"Ӧ:�u.*dg?ŝ<d[s�d V�E��J8nx�4�,aoڿ�z;�Ǥ!<J�'��A۽�0��n���
��$5�Ook��1��&Һ��<O(Z���Yt�i}�5H���t����-OV^�w\|ymF�a�e��4&�F�~�v���| iV�8*�Le�*�v�5<X�V���-`b�͓u�����Kp��E�l�v/��CQ�ٮ��L���L�}|smB90IS:�x��$�ɑo�y$lwU���^��&j�q�$|ȃ�f�N{�L�uJ��ޱ(�3ˀe�$�ck�&ˑ�ٖδqh^�"d$|��4,Lm�#��b�wJ������p+~�.
>~���d�?�Ŵպ���A�S	��#4�r\�3�ZNA�|=q;��&��h��{�]{C��i\|���ݐ}%�αx
���n���lC�0֊��e�س�����T���H�,��
1�Y����e�c�گ#��u,_W�67����'��@����+����-��%^��eF?�*C@��ɪF�3��*T�.��φ٦v3�[�?p�[њ�Æ����^��2gDG�.��c$X,�ƅ��:5�k仇޹l��{�%�3���i�>8�$�����Dv��B���VJPh�'�S(���*xJPϖ�k��I����h��|�OV�"��L2ۊv�*�M{�4��7A`W���5��k@H`>}486�D���M�	�GIJm��~"k�u6����a���ay��?)�����
2�pg~��>�?p���,v�-$��2>y�MBA����R`z�P�q�h^�/.����<)������|^qxr�y����drR��i���f(�~/x�V?%��=�W*��:VL��@����N�d8A���L#��χr)�pyvM`��o.�rf�0�������Ҕ f�����H���$��+�"T=��.,�Zd���k)�%J�Ǖ
�B�(�ӪPO-�\n̏����CRs8�_ɟ��2�?n7�&�Y�Vm-��ϣ2V��(h��P�
s�<�����}{��%o��(�%��'V��Se���d��@�����8���*U(	�c%�^z�ya��2�^Y> �j�u�jѧ�$����ruF�5�������<Z"U��,[~���o0�1ʪl<�?�e>��8�m�NO+��R<~�d^�I���~�����^=��Sȯ�� �s�]oSU��Տ�q^�m��(!� 8sNN�e���ܜB���ܳ���S
��c-a'wF	���+���<0��ZE*O�z,���8�-�0u���f3C�*;x_��'�8��WQ�z�����U�i7oqv�[��,�է�{L�ܡ���DrH�#?&���Ա����D�u�!�,3�r̳�"!�SkF$�g��"E�DV0je���]T�_ĐX�
~�ڢxd��6U���HIg�O����G*5O*'	-���gl�Eth ^�K�����
�g���8 �˖�5|�"]��9�p��X�[�H���L�n�-[�:�+�ӷ�^�_rC��F5� ���^��G7�W,8�63��MBY5�7S�<�Q�A*��TO(Գ%by����粭v�'�a+���>ߏ}�}����ɳ
N#A�O�Y��'g��#!m�%
ܑ���`�TB� f���^�4�W�_�O���2���ZIe�2�[?�����'�(�DX�!��G�k�8;wda������]u[�_Zb����̤D�:��X(�Q�kcQhS�~����3���O0��pwDXٲ�[ ���{b�G	�6�3 9b�e�#�������ݯeM�ۼM�K �O���x�D@��J�B���J@��dm��C�X����Yƌ�O��~�ڽ��+�u���0 '�1�U���{s�SA�����n��;���>?�L0�%������Is�$t�˾Ok�� �ڮ�*$Z'�?���ݮ���.����l��P�T�͓\�Y������W,�Pc.w8���*Ux~��ڱ��dd�Rd8�_�=��P�-#����WP��H��G�ث�y���L6�!��de��|8���9���G�����:^w)�\�?,L���kV� ���PQ>�c���>d�	eu���}[ZB=͛�]}��֭
��M�	"�<mXB �����O�f u{���
��6�[衮U�7�n��/d����	��*�8����Y�)nw��)ۀ�ٝϵ�>+��~��߰v�a�|ʞ���������"����|�ha�S���?\���}��~�<zٗd��{s>�U^�E��3�s ����,{�#_\8��dk]go܄��a����3#���e�a�<�����}�d��Ϭt�	�P����0�W��.�qe*��.�J��Z�ˆ�枣�i���	�����M}3�@����B�48���{S�vl�.�
Kov��-�':��蜁����"�8���zv+h�6-4@�߰����1:_ŀ�
�nqü�f �}V:�q���]r��:�쁒P Ժ��Y3?�]@��ӵA>5�mm����]+��W��!����|��W�n�ܔ7����#PK:6Q��/B^��kz����S	,3�f����T��l���i��="[��-��4�:L&�rb;��$ᜢE\V�n�'��/�0�!�r	��ob�zÓ����g}���/��Q�Q�RcovWG����a����@�Up[=Zê��
��u�A�i��6�X�C��x{?i�$�D�s���,u���6�huZ�
9�����5Ϗ	ӑ�E|��چ1~g�st�ˆ���!����a/���������L�/���.	R�E��*ݒ^Rd=Ѽ~�ghma����,91t;��\�>N~�n�YA���&il�,n�v���R��ϿnT�w�Y<�/�������?6��5��S�d���"��1���4�I�8�S�E-�p�SyT���H�Z��W���(��ۙ,��7כ�֙��.��:N��kC��C�p�'2M�T"�}ԁ�"e5�]�;&�MiB��.o��I9饽�,���&m;�g]G�t{C8����[w}$^�k���侰z�(�������X�`�C��`��j�ʏ ��O��VJ6�@s���M6i�3�5��"z�=���9�e�Z�P���r���P��]�+׊>z���c=P쏛��c�})u�������C&5R�ڼV�PQ�N�����3ԉ����6����G2(�l&�s���������[�l���w��2�[��H+؄�A�U��]���;+vU��)bGy�����ޜ���:���� ��4�ä>�u?ڞ����-���:����ޫ�k{퉺W	W����{�.�ϓQ�U�>�D�à�Qq�j����g��nx_��ci�ݙ�I?���`���pF� �������犓U�19U�Zӽ�uJz����[H�u���3���N�88���!&�ůr�p���d Xz��!m�j�p�]���r�|~sSwvX3�x���
n�tJ�跖��x�t�82�=zE|�%(�@�O��d����WoR}�K�݀�������A-ϔ���$R��9T�z�B�rG�0_j'�pa"�倉�7ȹD�@XO��.K�5�����~�pTAj�'�_�s�~��A�}Y� mh_�/Ɍ6 �=h�b%	Ɇk���E��q'�il�}T"Y�p{�k��t����;m�>M�z�'�-�Z&�f?u';<�M+���<1�q�����
��4���q�m���i��WK����B
�l�ԑe1�w(@jZ���9���ξ9�\2���\�FN?��
܊������?��`�A	�i��ځ����,���Uu�Oy��ql����)Y4�wK����=��^E:�1�>P����x8?ZX5�^���4��W8�U��4�ډ���H�$?�&���S�����9`�ON��=�p�݊ ��ޭ��`�����콩��������Z<��&2�g7_
^7�ߕ�>��"�^t`�x/e?��t�q���� �x".*y�C{�Z퍪KpB�Ex�C0��F��3|pz��R�=T$��uvZ�U�������} w�ҟ�����0�u��a��~��<��]�A�9��{���Yk���V����A��*#���%lʤ���B���6�]�!�:-�X �̇t�&P������~��#T�r��$x;�D��	��5������n'￿�&��V���$D��	CMp����b�`����^Ӣva2w�]P%�S�wQ�|A�&A^h�V-�M^ ��B������?���qLҕoV�������)�c�*��������D�g��n��l�0I�0�$�����E���tA��7o�n's��j7Og��A�Uo�&I�Z&�o�Ӕ��%� �e>q^����wr�m��c��/k#ݨ�5Je��٣�'|-A���
��60��` ��|�b�H''�9�|T���n��σ�/xCV�%�({�����\���-Ҫ�T5DՇ��ն�'�f�������=��a�L��?��RU-P�*r��n�+4�zQ:�M���x�>�>�����D�aI�ߗ���N�O��㾆��?�7�:-�9�::�L\��p�7�ֺ����X�u?b����p��O/;y$gkW=Y�K���#���"G[x0~,
�<����S}y ʬ��Ϥ��+_w��8f��2�L��AKj�9��<�B|v`�P�n���.y%pCT5�O<NS}��@�|!ǘf�z��G��G-:��la�?Z���r:�9z���!��4F�벬=u7˴���gemOX�8ǧ��בM�=�z�Z���=Aϣ%{�J֮�Q?43��Z�eF�`���mE��D�R9���[�p�6�q�b9�7��ma[��o�ǚ�׈q�ű(�]1���C�8.��/�u�d�
0��S�����͗����x��x�Z�����<um��w�����Ȭ�-�C3=Mi��cW�Wp�8�CF�Ҝ��[��φ:�����_\dTV��?-;}��{@�������0%㝦hɲ�[2 ��#��6��=�C���X4���^N1�pc=]���>
�C�����{�6�k�8�vI�5O,�1S�B�~��0�#�5�F�Fg]M���R�{�h�8K��H���ГӶW�c�7ڷ�����߮��2��3�D���l���3ƌ�bn��ܟv���aܽ�����a����`�z��dE�x����U
ɽ����1��u^��mo���"��܏��-���9C�ij��(��-�"�K=�ҽ���y�R5N_(vvi�*��j¯uA�k��h[{_�g���J�w�g���>B>'���N:��`�*�zR�D��4m�[w��¦߬����<\�eެ��rst����?"�������1��o�_�K�DT�4��a}h�`H�O��6���Nf��u �%�ߕܵ(����f�	���J��L�q�nzq?Bu����uڻT�6~���{D8�#۽�&��%^&��p�VX��<8��0IcN�Cc��B7��Kk������2�lr� C'ym.k�(S�B�%����E�Ԗ��l��h��R٤��ș��p�u�]�n��<��<j�ҊU�N{�^-�5T���Ź*�P���w�]G�������z�7�5;�~��sia{Q'_U��~q\y1����K�-��2���D�o�p�?������n]-����W1��@RX�wS��1ɀ�T��x�f\D8��.s�&$߬ )��ȓ��.k�aK֩�hё{n����h��bN���oMr܇���,�,�XNCT�p_�k}����Uɬʡ�k�̊��L"�ח�>�i�4f�����l����<[���e��w)�+|��s6#/Uq���V:������%���83~f%,[Q��R<��ې�&	9��T�Ƣ�%] L9�秌VMU�.P���>��,�Ζ��d�WC5G�7�Zţ
mli�waM"E�m��8˹8���'yf7g��6ZP Gxt�z?�ְ��y�2O��kko�io��4 f�}S�V81A��^�����:��4���yP�|�HA4^�����'n����7H[�E���O�Qju�Qg�r��齱;^��z��˞ɷXj"z|zq|w�I�V��z��CB~�節�;+I��96�b��J#����q�F&��eY�q��h���}�'4g�2����礣<7H㫳~UI�+~�*��m�쎗iq{h��)��Gn
��]"�!����Ԧy�o<��ӕ�ۣO4\&3_�
�VE����*�����>2ߢ����.����0Re�@�y��F��ۑ❭��ܣ�s��\��76Hk����¨j�P�6,s�h1�3{(\�n6�v^�k��}��A杓|"�"��]�AI�	���l͗^ͼP���M��C���p"-]�D����F�)%��8B6��!�%��]Ϝ��8����E�;���j�m�2MI�/���{��,��B�Ƙ�&��)�(�^ΚK^^Y��_�#,us{|�]4�|��)U<� �Kj~%��IF��4�t [��2��VE���(��Yv��~�|��u�I-ipr��ԧ�w6�Y#�[qbfjyr�����в�+*�#*QǢߺn�\t!ץ��u��/��W`!�l�n?�ʬ�GÁ�����k����ZuA�ʳ��@Ȟ�k��K�\F�ڐ�|d{�Ⱦ��3|P�2Z��YqP=#SZ��Gg�{�����_��҄JB+����=�n8靧V�5�v��Lu9󖿑���� ���!���gWw�l��abPS*����k����_2�6���Tg��Ɛ��q��̱�J�ş�Uݓ�{�h��Mx7��4΋{i�fFz�ǚ�1lh�S3��Y��e�A���=U�E-��Y�����
Sj��;��0�cCǷ��kD��<UB���{{W�\���Z��;�I��r}P�grʊV���8�k��6N���wי���\��׋��wf�����\~dK�]�5V����|�_�G:NW��B{��?��6��d��ڊ�.�槚�Q�������v�䈪�s���B�O ��gz�'���*=}կ�!���m��8?;D�7<��>�']!�����U?5.OQR`��>�_L�>3�R����
.�o񘑘�=B�WE/�x�:���v���7^�<�M�����@�u�-B:��K����A^��ff���, mx~��ۿ�x��������C������
�o�# �e����K
؂�%c_�Y1�+3w�	��B�&go�J�gLo�6)�`gC������a'b���x�E{�?]5��3�Y�QRp�����J������a0r�����xPpyg��dsy�.G�^�?�F˅��S�?� ��|ZN����z���U4�p���F���'����o[)�����p� �l��j�;�+���P	�q��+p����߇I(Ar��%0��YH�mQÌ��T��ΨㆸΨ�o����;���Q�� ����r2 `�r�c�����q����P�K�s�I����V�ݘ�|��;o�kh��K�9��x��񰯦���s�_现���n�C�DO���B���ԟ�^S!O�n�N̰ho�O��6�I����h�\f�;,Gw����B���>�.���2_6��UHӬ��.ֹ���Omi�����̾`z�ed�8)��]�l;s��Q���3 �.(�����]z�:��@ݝ�������
�q"���[Z���fo,����/��.E.z�=ˁw�7��S�7���-����j�����DQ��1���iIkW�L�4�P�sp�5˩��"/��Uv����o��\�99��,�������i��FK�Wx#�9�AGVV.(W/�+7ڻ��l%T�	�(��NBL�C��xЋ�j��yL\�p[Uj��.F!��?��jʢi�^�#��*�$� v����'ۛYN�VF���~����4Btx/v��J��������r'�d3�طb���e�dK%��Cw��Y��2�<LNY��b3�4��֒U���S�*��g�-,�Fi@#��l��%����JԷ�_��Uգ���)�d�wr*�5�5I.*�p-ӓ��Ǭ��Σ	��R�]�I]?���MW�ؗ�,�ɬc
C7c�����&�	X���l�u��k��6��|<{�^��d"RItf�-�X;i����'��'6���G{xꊲ��p����"�[�����N,�� �]���O��
��q�z~�ÜN'o�/5ԩ���Ǘ��P�%�{��/���X�b�T><�/�~��=s �5�c!�B�O�L��f�aS������`+x���vf�<��[98������GW���6Nm$�.�-<�Pe�V485�W�o��(�<?=w�|�h߱��œ,�c?����|2;fｋ!��)F�A�N����	u�O�j��A����'Qi��i1�ߦ�%�v���A��"?�	`�JOx��ҏbQ���g���2�"�u�f'�m*���2�)k���6f�H�/܉@����ԛ�ܻ�ʌ
K޺���S?~b��n��f���;4�H��o%/��*���k�QT��/u���v3���p����r]�a9�1�cB�]���zu��	ޫIF�©#2�(���R���r�)Ԗͷ��:��}��cy���Y�)q(+��+��Y���[dȴ%�,Z�~���u���[���R4
D�xy�+�|���?��f��Ĥ���/Q4�i�=z|�7��*/���.���ug��Z6��CЃUM�xݟ��oA_R�u������M�� 2�mW�z�,
��k��5�1��?�����J�n���ڂ�W{�k�ž��}/�n�']Ԣ9���۵�l�p�*����#C!_�qoiw���TpB0�)�ٹѫ$�s>�#7e�}�ڷ�f���$��������W8l70��e)�ß~|��1��N�����$G�ܽ���+Tk!3�!~����'{��"n�,!�W���h�<���ސ,��M�@o���0���:�j��&7! �$R�ke�ͽ�@���!�H��r�ݿ���h�-_��-�j�)pվ�*F֊p�F�`u�v�$?��m[��~ٜE�RB;N�D#�F�@�;���i[�Jӽ��5��oG��ĞykV�L�����|A|�}�7��fb<�o��vG
Gڨ}E�0uY��C�88��jCHO3���ſg�a���}[�����n����۲�SɎ16g[���$˅�;c�y��0��Y��X�GDkA�\Y4�Z�Y����B�W;���*��Q'*�F�w��=�ϔͯ�5�O�p�4lF%�b�e~���T�H����8c�䎲R��܉����^3�����^vk>������;;�x����+iOa�f.|t�H����S��ytˇn��E	�����M����Ux>H|(�O�P&w�0xW7��Aȯ%���akm%��:��ʻ�0��7���5ot��(ܥ�����R��Z�/5�̄�^��A{R�F���d���t�$h�i������ݜ���p��k�56�n����~��Z:ߋr�%�S�m��ClO�w����N()h�#7p�V�4Dk���/�Q��C� )��_��ـ�����b�\�E���l 鏙dDA�E��J�<�*�5���C��;
�"��2��¢Oq�K�{��3{�X�y�.P���������~L��*�E%��Pi�o?����h8��u)~�b6z����,M��]�Ÿy��흙�H�7 vEV��6��uE9��y�.��=�9"A+�}R�<P���ď�sSqy�����X*=K�������ɺmP�:���o��s���s��0_RIf������^�d'�}I�8M��Ne9L�T�k-"�;Aɲ:��d��W�|8j`P�S%Σ�	�qK����/��bv�A��
�J➣�d򑿍�)��*fU E�&��Jn,:��-Ol����=
��mgx5���ě�4iȲ�JC��?6�wΚ�c��k+�D_�g�t�����n�&�-o
ͻ+�����w�2d�0�aà�c�Oܮ���F�U�o_���?C�����:�Ӝ[�;)P!�W`���u���� �I�`u4_�ڰ�t�l�ȯ��6��<�R� B3�h����!����U� �x�?1��qȭ;:�Tн�IV��Ԝ����['�����tU��?���becs�0_���{��Wf8��'o�LB�7W���?T�)�is��'��v����xB��شxu�-��]��S��Β�W�`�b{w��	��Wx���^p�4�4��$��2b�ܱt�l7S%� ��+B���N٥���ȡc/�A)�Ydc�,��"����q�ç"���&��X��M��̚��a�m�;IWK�ixO��&-��8�ϊ�DD���P���m:`�3��ғ�t��@[7\4�a���B��O"=N="�D��Em��r���F�m�ڱ���+�R�t���4�ԓ
�@�N�ܮ'�=y�������?D���hv����w���*^��l��BQ��ְ����s��F��%�x�eX�R�lڇB5L���g��n�jF2���:�2LFKyJ����7m1n��
w�k�D�8�DȾ�5|�z屹����?#���]8��(�#U�9/���K�R��bY(n�����Ter�9Q&Xn����pk�lk����bHd�C�}8��c�mrvk�l�0dL�&���ʗ�:��i��?�{m2�G�F/F���z?��gƱ��-l��ݥ����~{?��7U��D��W��꼮6���)�$��&�)�����Vq�.����3.�K�k�̩%$R����J���x ?Ie��\������~l��$%�&�R'��l�9[�L�6&�� ҃�Q��{bl��X��X&�i���#k2��e";2	xzl�8����֩j4U�@��(Z�����4tnA�M���[u,�ŋ}���9�^G$Jː�kϪ����{�� �:�6�����qvś���7!�c��{���[!�G��}�	�O�������n�_TA?� ��w���?�?%%�ރN��M��2��	t�i���	����f�vX�����W0x#y�O�u:T3�ۙP�
U��\_����l$���#���x���i��ka��iQ�p�&������O�'v��I�Wn��"5�|ӿ���tȫ���M����o��U@?��jݷJו��[]�H�P�U$`.�m�lB�#��f�be2�}���z^ ;������&��\*�][�ъ�ֽ�zi��Oֺ+27�N��C���A�W����c��Zbd"�ȭ����n~"S��[R̽o�!8�b�\�� �	��j��P�~E9v��54)�ciy�a�*+���+N�k�˓sߝ+>��K�����l��t^K�h\{7���/-Yl�G��0Q�����D&zj�.I&�|Ȍ��&_s��ݞ��4 ޴��
_h��,�����}V(r�ڔ[�>`��蔆���A>zk���0n�_(�ْ�m�Q�q{���Eof��g�t�Ը����oe̓�>��UAC^�27�҂Ŧ�oȰ�h�|�{f[�H�=yx�j[[TkY�=�-�X˗�IR��ѫ�Y�[T]#<�"��>��H������W�� ���\{j���kΈ-��c1 �SX����+\��FE̜�ǻ�~=���t
L/�w�gaW�v�Ce4��A�S����W�������3=e���ˇ����y���Q�8�W��/��P���'��c Q�lQ�o�D���ψ`x��_�!�@jWC�W�y���Aщ�g�<#Ҹ�t"VW7Z�	�΁��蠖�����2Z���H��H�Cw��Mo��f�n^R]A����v�����.��F@��fU�~ٚ�,��V���`��������rV�ԑ  �{�'��i�\���W�!-<���0�O��v*�����g1�kIɆ ��� 4UȖ��u�~�5fL��y��i�2��p��{J��פ���������hH��0�2c��[el]�b�x.Ư_N~>-pP��ƕ����[N�Y���"��-�*�VC�O:b�^'E6�7���9�J��*�z������`;��5v�Mgj�����lk�2<-%����i�Or�������Wg�M�r�����"�B����H���i �Nh�����!V���	㴆8̐���⌤�־�G59�JK�3���;�4�2jc���YÐr��2���R��n�����R%���E�Ǒ9�X���aYd��b�?�`A��^��0[�ǈ�a�6.I���eGѫ�M���5��W"�&�Y7�ήl��K��A�]���E2��2d�Y����3ZI#oPE�F`���#x�%�Խ!���E��4�V/�Tfބ�G�a��٥���m�p�S�h)�Im#Cz�2�C�*�"�M}A!����;�Q��o�8��޶0�(��+��>�l�Oئ4h��ʻ�� [)i\[:'���m�l�u�xQ�����#bqBS&qq�پ�W�u}��
/_\A.��_մ!M�bn|��f�����u���~���ĲT�I�������7��Q�}�v)3*K�&�5�ކ|��;���X)��k�-����3���m0�d,�uW٫0�)���!��hF���c͋����v"�>��P�v�GN��dq�6� �5xCr�7T�,k�HD�b����3������I�^k�����DztA��.���C��^>��V����:�(&�f��o��q��{��A���g�a�/M9K���|�"Y�#"���`�� �����Ozy�GZ�޿=!�����)|�X�1��2<
�_۪�EV�<s�������i#�� R����t�|��0o���s�0#�=�b
�{��E�s��6f�aa�9��l�-���:U�1��,jZ�à��������뚍7d1?������^f�'��_�G�C�_}�.{�Н�_M#I�8����]q�ՓYI8�r	(�č#Bn�*Eq�s�Zhn&���њE��-��t˕�D���e���vv�Nyh�?U������Sd���[;cΉν�zI�>~;I��M֛f����V?�'��Ui��7=�&��V��3d�N���]W�?��� Fǎ����Ѱ��Owc
���0�_j�?]%��b��2�ц��(-+�Mb���m���m������zH��ӓ�X6t�~rA���*���5�����LLĥ�_��}E#S���Q�l���`��8bS�H;`�j�[A<e�ZsP��8�W� <M�s�-�^�r�7;?�k,�A�pp����.F��R&��H[Ӭ�vk:n�Ʉ�}1��G�v=D�*�]��)G�Kn���(&>7��o�2A����'����CpXn~V�q{Wf#HX	ޡ����K.6+	�P�X��Jeބ�K�a.PZ�$�܂/ki��AIa��&�ݣ�!��4�[\M���%�;'�����3��4���C�dpw���·�����]u�=��W��Æ�#��A�>sq~�5��o�+��j�xkL�cA�a词�4��A�Y����:�3l(2E��@���{"J�#Ah�i�:0�S?��H���� L!Y��:�F�U|��pG���Va�eJQ�'7��7�������7Z��S�e)�_Ң����f��Y/,�Dѻ�I�V�=~�%TɸV	�������3����R���C�[��"$�ٌ6�v�X�@��ݟ�ek�##�gZ��.���q�5������ ���*���_�)�>Yǐ��C�.�#m��n��!"�9���ə�fA�������e�#�Kz�K��N S�0�XD�U�#���Q߆�UT>}�m��*��t��q3ej��K^d��IM>��Z�b�z|�h{��:"칡�u?�p�x�G&���}�k�G�{�v�!eE`
dJLȎ1�g�RT̀Z�,��)3�3*h�Ei��u=�=�M�~o�;̮�V̇�X��-�P=n�"j�d���n�G�i*�σ��;W
eeU�������Tg��K���YF#~����Cb�ŷ�@�!�FC��o��d�?\'M��ۉ�;N�!r�&!���&�<Z�v���B}�#
�9��@�H��\��ձ@�S��WRD���<���]�����K쓾�X��KԌ���3��k��n:���S1��O?�����s���3����F���5&QU�=���l�O�(Ȏe,Fm�ҡT�c����^�c��i(��6P��`<�P:�����( cĴ4�*�ʓ�灨X\��̑�{�Ҳ�'W��$&����:Fk������D"���Tۼ�w�Hr��Y���Sf����
d����}sbB+HT���*8ʩ����{�Z���U� ���wŗ���I]�p]��+������d�4������XQd~��:@�K˩m��?�8�%j3����þ���uB�V����g�}���37m��'�4{hD��/���ξ��'%GF]�������O����G�hH�v[���G������ea�b���tCR���:�N���)��_�L@S�H��y��Ǐ+>�P޻�(_0������w�u����娴���q�1��Y��@�3�²�A�V�C�7/�X=��c?���D�.T~wF�$K�Z�w#���x��t=���`�G�h�k�#�i������ 6w:\N����w�)!X�^��
p�	�M���I��eڎ��{��p9IMg���֬A��@c���k�=[h|޾^�4��8�Y�#q�9.��
�%��!�1�V��������M���b�ߛ
n����U�Uydw�u�� ��ʷ��t���;ΉJ�m"�M6��i�G�����FW>�w~�c����ϰ얊���<���is�h�P�Ǥ��9�ٽ�����E�� L�4.�en
�ԧ�7�������
d��>)p\x�k�6�B�=u-�Y:�-�Ur���yW���̬>oϥ�BV���*DE��zy��B�
�Di]��U �`���%o�Fg�L���kL)%Li�����������2�����>E��A�bT&�Z��KA��%�Bwd�r_e<%j$ƀ+����ί�h>�=ّH?g�o���Yˍ�_��[����x�!���e��R?��h�E{9��.�P��jY̥��.��-���n�r�I栊R���Pk(9F�w|��-@h��Gb����|8�{=��Ю#�b���ڼc�#%]��))�� ��Qp,�K��m^<au������[�C�_G�����jr��zm5�����l������X�f�ey�>F�GRMj$�n|�q�H�B�m^����S����ju^��`$2j�[U��Y�~���v�����zB$�"|$+���� "�{���FCA���#��l�����,܎��X�l�6%�y�7��3\lܩ�~�)���G+�-�x�;���g^
�A�-�h!�F��[��0'��/��覽��,���Q/�T�w����ug��<X�󎼲Fe����]Mtd"AE��>8l���[��-�+)�h�]S[r� &T\��u�,��L�Iw'�ʲ���#f����O�P5ٮ�2G���3���C�,2��j���J�����n c^4�o�ї��d��e� �|KIֽp}e�gX�K�L�״N<D�
;�h0�zc��l�H��2��QpԾ�0��|g��}oN-��+\���}?�qQ������(cBBU�?6���n��8m>y�}��&�������C%�.o�Za�Q,��o\��-�e��Ә*���t.��͡RJ6���DEjL�KS��+���5s��.V�'��P��_���|[���<>�F�?��.�	������[��g��t�%�z�>vK#�8��}>l+�2>�	J��S�kP���F�G�kˍى�\؄�	m�;&{l1���o���^M
78_6g�Z���z~ �;����֥����f���kF�O�FZ	G�!H�m�@&�)����cN��Z"�4�^��05�q�����2b�����翲/�`����޸/P���ǻ?b��̚��:6/����N���^Q9�S�Ch_�<v��ID�t����w�x��JK��)N+�9 Yr���B��o;!DHb	�����r�=F̂c�,ʆ�T��7�%^HpphM<�����Cm@D��8���.�?4�q��ff/�m��ib��Sc�'ڒ|�
��Qew���xj /o[�/�A�>����S��m��R��.�xx�a�#Z!Nn�!�N�58���6�lU%����C0��-���X���%I84.�LY�v\ޞnѩ�;X� ��.��h�
���u�B�ڦ�;���<b7RM:���Ȭ�+o���t�`Yr�U��3y=�{�������S�!v6�N<��_X�����j��,l2D����X�5#�Ȭrz�w}#x@�;'�k���#�7�/>������G�����\3�n�fy���b��.�i)� ߐ[� O��/��ꚗy����e5�uU��Y�Z�Z�.��U)�@4e�eA���LT���!�[���<��v�	f���B֨�`R���F�;�D+b��f�nD������Ğl>oV�������L�&�/�����v��86׭&AL�b� �asdb�L,uɲ�4�z��8*GH/���f.���n�T>��DN:��$���uV�V��W�$K@�� ��<d^G׈6��3�x&(�X:a9��ܒ�t�������Z����*Pޝ������n�;u!x��9~�d/s]���O���E�5�c[�{��A엔O��h��V���ׄ[�l�Qܕ�id
ޥ/l�H���2~��f�H�<g�b�< -
�!h�rO(0.�+cP�(\�ź�w�i���[�����6/J{H{�dk�4�j�܋ۯ�<j���X�<��������k�D��%
�1s�p�L:��YN-!7s�+�o�hiÁ�J+ ��<d�)����ްI6�q�Η	�����?�lg�d��Z�Y�7�E~̝n�߸��kXm}e1�i��K�'�m��|�n�N0���ݮ��\O�帖�Hn�~��\�A_�&�+��N�����!h\��%���Gg�T�l��jx�7=�e��a���@�jdI��j�pD+��Q(�%	E��#u춣 �
�H�H�Cn&����TM8�H���c��-?@�e�{mٍ=��p»Z�Ɣe�B�Mb}!�����c-�>��%؞	:y.�l�u�U��}�a�Z;H��c:�&/�*��;�S�/!���`�NAifb�,,6]�"hq/p���� �L�A��Xÿd���}ƕ,A�%n7C�*$������I�<���͡eTޭ�Z!�t#���y:�ƞ�y���FZ8;~�q�h#�:�\�FE����<���:5Z%�RIO��܁%�sWK��.��]]ś\��Y���\k���z�:,�U#�N{��!E5	�.14� a���p�Yi���|I��lx�m��6�� R�����]�`'3+��侷�����y�����UN�`[)K�Arnl��,I6��d�mq����KN�☠�����y�3>m϶N�;J�7�	b1��pv�|K#t/��4|�`��#���}RG�94j�boO��LM]@`�Hrw�{��%?�����J����!��K��uJ���[���*iL�7�3�/�F�8�-Y�_sP��Y���KӴb�3a���=�<;��Q&r����䩳�5d�&�����#j��c��8	�72��˭�=��]^?�ݎGԳ�;%ѽ��bh���8u��E��!��}Ys
�8_�3ٓ���h��#F��N�+���"�'�6���h�K��k3����(�8��T�)&�y7J
�Ilx�ԶR�5Gu1��e���~ɭ��$
}�÷(�)2f�`Y�٫E��#4�}C�u�K�KD�Ma�O���ְ,�<�K�:Y�l�m�$�6"��0#�N�"�'I@�j���U26hZ��'�}CSt�1�1�nR�;��3��/����J��/ى|�[�?q�$Կ�2�U����i�J�3D����r��r޻̶�>i$�0%����j;6�$���I���K�����ތ��G>~�;�o� ���M�
��qw��m껼�L�X}g�e�p����6(Z��U��BGS(�,��8��R{�L{Y�?�|9�ҧY7��U�X�4ɠ�$�f���p&���o��!g��Lͼ�_7I�b`<7�C��~�N;��t^�7�4I(���\�T��\!�4���G&�K�&�#,k	v\��s����FNm��8QƧp/��+�A� �1���ƹ�~wa�v�2"���`���6z��c�6<�*O� �[��p��i���Za��.��Гߘ������� 	a-����]-�gh�7�]V�7Q���/��u����ysO8�\��-���n�$oeBe%�B5ͤ�zXLe־�s�M2�	�x8�^������v�{l&v�X9Rs��L���r�f#�Uv��ʸ����ߚ׭��h�3���u���<{\ᘩ�	W>����]��X\�
A<�-�Xam���*9a�*�C_o@#��6Ω-����(��I��	�a�9�����w�����=-`竨'݋;fS��oak}/�'{@>�'|u/����ɑ:���9,X���5�^rrp���K�~��%�#���-���7�E��7{Z�uH�Uj�=����f��X�05=����]}�>�P�{�D�7K��E�pQIW�F�Ϋ�zh�d�'���Ϯ|��&�����v�$/$2�f��ܼՁטq:L�9o�]�c(�1�E�gI��J�e�DB��#����\���)c��2���I2^��Y�-�=���O����g���ҞK�U&��箄�������bBO���^}��y5�M��eQ+4V�IO���^�/>oKc���%N[ˣ>�|�\���.�im�-�sNݬhy������`�K"-A���Z�2����_~^�E�w˽  "UbTb���c�E�]��z�S����H�A=��LSO��{�,˥;�#\Lk�D�z��=EE���"��x���6J�[�=���Pό�X ]n�3)�'���74�q����&RXp����=�G��AFK;�k;�8G#��w�^O�Y�-!�i;�G�4Y���⤉[�?w }i��T%Y7�]�RY�	yǾ�M��X:R6>��e�Ug���W���m��Ze�!mԙ�&@�o��*;�JC_����x��ն(�wƲ~d�I!�� 4�[SO�J؂�8}F)�}
(f vq����|Wi�����e�umEbИ���\z�iȸ�9�m4�V3�0���R32�^E��הK�����5�p'}��A#�
�R�zD��Ŵ�b`X����
��)Qi�#���q˅F9(:��<�ERLXQ9c{=%���@�#���S��!��g���>~�+%�mB�.1%=�������M�X6�"X?��4ظ}�Y8H#���g��Vr��u��ॅ��H��8iS�Z!�`}K|��������)Kww���!Ο��)bu��93�	��^�=28��f����
g�,�7� oI���ة��8%;���R:������� ���g��G�7?�^�L�,gG�֏\��T�հv�=uN"ZB�������".�*O>'�c�9�8�z��g�jN� 3	ALdZ�om�K���zNr�Z�i�Y��|�w+��T�����&�+��V�(�OJ3���am��1���)K�o�Z����[}Zz�z�������gw���@m�_�
%�K[+��q�s�� ��:��|K�$�'�9Wx�4�������Ӊ[ܴɠsU��T��v���516"SƯ��(�C��B�x���t�R�T��o��cB�N�۠���)�7�J4���h�K��&����J�TvR�(<��v�5�᭢e9N��%�tX���e�G�}�����u���?�c>�������sn��
��1�^��6_ށ�ǈ�@�%�l(�c�p�bk�7��/emx���[M �=�����#���ȲcZ����.��İ��3�v���W��r0k��C�J�����n�:��_�"�>>���+Ү1P���P�{���
�^�5���ܘ�����e��*��}X�N��<����{����+�y��h�x���+K�O]t�.���E��w��[	:9\n�����)a�����[�#4/���j�kh�c��b�1+�s/�6Ú���߭,3�~��χ����9
;��F���)��Q�u �A?Ty���T�c��w˭��b��D��vX�3�|X!�[2�t��'����d�@�3��%�QD�uM��V�e�h�7π���j	�1�Êm��_ � ?����F3R�O����3W@�Ep9��Ca%w�{�p8a_5	�Ѝ�e
?�v�W�,!Y(���_�'V�Qd2\${�d.K�q~��yQ4/�]���Zs�4���[���3t�}�Lu
Y.�m|�_<Ny�p�&���9���s�Ȟ�;H?S���HB��_��l��� ujz�ƾeT�6^��ܷ�	橿wdg���^9����6�M�f"�EիJ�q'��}vaY��P���X��)�M���Q�["ݡ��e�F{}����F"���ȴ���:		�(�cZz=I)�d t��X��?�ʼQL��D?�ylQ�fQ�{\G�)��c~�:: �	�K��V;�ȏ���\	����ѧ~>��E��5ߋ2�>��𢲻�p��V��:������3�~�����f��#L1h�&��Ȭ�����?Xh�5�xt�]%0�tIP9�մy��o[�mV!j��ȟ�U)�M�g�f T����X:�����-F+�G�m�ͧK[��6B�~D����x�|����;��0N��t���湱��Ǝ��=(NVnz܆�����y;�����a	�|>�1̸���,�)u���TU0���ɏ���N�����]О2�su��-�G����v}X�{�Kޢ��w7'��p��]>l��\��C�4��p�z�V��h!�.Y�ǝȣ����[쏅��cXK�7�P���H�}]fA���d>M�'�΃��֤C��8l��&�Ӫ[%��>#zx��u��8���h� .~��8|���1:=)�+�����9}�C��]�v�JW÷�KY0l���>��A�AX\�����{�d���}���Q�r���?���T*����(��A���K]��*Zr�yW���/xza�S��H���VM�o�����U�Z՜%�8�9O2�Q�����U!xy�D$����suNk\6��IJs�����Q��lK�G�b"�_���B��YiU �=��S�䮼��=Zʻ�"a���oA� )B]�a�.�
_u���_ڊ
����X���ۺg���{c=H?M�/a
ML����G����p��݇U�R$4�3�,S5�*B���'��)����
�/�pd|j�4�A�#8�.|X�2��O�Ʊ�K�NK�_�_s�o������&"���U+�.��|�Ge5v��w���w@��7�K+=�$��̕���
Gp�	!`�E���ǥ5م8��fD,-8,G��DC@m��D�/L?�Lع+T�#��U�1���d���6������{k'�~&"�6�=vC��ٹL��"vq�9۟rׄ��&�|�),h�e�2L�6LW��gU�dǶ%�4J5�2Q��(:N�c)�f�W���|���'�O�&ߦ]bJ�=1&�Pۤ�h�����g��h݆k&�G�/vb�ڜvEi���(o���)�9;ݻ��AM��OE�E�.|�%u��� �ҥ852��ж×bh�����A�����%*7�T}�K��]4��?+��X��}���D���Z�B����c�g���M�R�s����	w�pr����ݴhֹ�?��j�]��o����w� ��L�o��蘑e���/9L�5��V� ݝP2���F�	X���M�����<p�Α��V��d�6KJ&��*�ڲ�`��eqW( n3k�q��,�}�{�O�L}H����ׇ�<~�R��1,+�R�;&f���h^��ߚ�m�M��ڎ]�p`����j�oo���z ߹�G���F�:li1)�v}��/���8����	K�B�������bɘ9���{��6Po�I�jh^��إ(O��g���`}���J�T�b-m�xS/�p*:J�s���_񫦂jqZq㊻���QzKv� ����t����+�kO�"�D����^@������e1%���s���ݶ.C��>�0V�o��?�8rȢVC��Ա���94�6�n�n�[�y�,�S��A/B�����֨2[�Ɓ�$#P�����,K��V_FB�B� G�G�j5K[9��\	X�X���Ŗ�^�P���p����
J�*9�榿�\s-
n����r7� �͠�����t��!�÷l�}u{��"��G��*�F2X}�}��s�g�E��_�"ujh�W�V4f��<Wg䥶���.������a�Ŷ�ñ(��]�0o�1<]�n��b�ɛ4�7���+ �T{4Dh�3�m��h>���;��Sc�H��~�`��%#-��Z����������Z$b������ͮ�L�$�/� <�^<�[ۙ ��/V�W�Zvw�w/��׵T����a:�2�G�P�1}��V���yb���~��?�t��[.yO���g�y=�"��4��Pަi�S=%��(���V/�~�%��/Cv*��#p�6��p�k�����M��޼�㤫#�,��\��	bozx��`�ո��o"�C�I�ߛ��TM����5��j?�D"z����z�ơHN� 6ҕM�Ɣ=Q���~ra	3�֦�N����W&���6Y���̓\����[���4�Dߗ �!*s�a)�s�cD�d�s���ո�� �@�5*ʃ>�{ƕ�B�ڥT��q�oѵd6pf�*���s��N_Ew��eB�f��~YԨ�B���}uu@x�`��zq�A�U�����I��,��������&�|�V��5Ą�e���F�����G������ի��Qgt����[2�C�m���ݖ%��
���a�M�6_��d)�'Ä3焵��O����[�od��-�\R�(S�}�����kS2���	�p�8:�[w�[��\I�c��r�I��>�e��eT4�g(�]*��݁�A�*���7~�&��M]"=1��"m�ط��5�V2Pa{O�6��V`W�q2xӀYI���i=�L��eג��sژϷ�qj`ͯ�a�3���æӜ�FW4]�E�+��,@�b0Z��"��knԈEՕU(o���m�_&�K��M�ki�����X�[�6e��ӕ�]�{�|9,Ȣ�s��gw�b�O#s�Η!��+�6�V��4������]�$\����DIX�~�o�:(D�:�e���J��Z��q�i�|:�a�>�!�fK�4���*�<���0�-L@P 5�ҝw;R~z�U���e����`��[l�)8.�$� �r����ԋ����<��^�e�n�u���O٤b�&�oɣ�d	K>C钙a�r��F��}F����Jm�����^A�� �yCk�
��U*h^v�G��_3#��)%⧌@lT$l�ߍ�t �&d�ک�G�:`i��A��c�o8_�;i��OQfq����Dl�g�L�Y������#�\��m����5d�t��]ǮSm��|:&�'?��U|�$��3��L�^���환�B�K�b�	�8�g0�N\���Z�t�S�BB�h���̞��1�M���p{�Q�	�"��s���Y��Cz;Q��2|��EP�gB��FW�a�&B	�Ȁ�bd�ˁyS�<�pvp�K�h5�ź������,�����cr�?�G��%_���Vo���+�380����A:Ș�V��;��*�\�E���s`��[6��}|��T��&b���`��A Bx5������c�E�o�m4�i���$��⑚����%��ᐠ���l����������'R���Дs����b� �I���f!.У��"�%����SBi���A���Y[5�Yv��O����u{R��q�߹P�&]�$�W�?%�?W�%�m�*�B����c'%q��tMqw��?���$����K��B��< �1p���J�1��xb�-5�ĤͰN& ������G�k�.q���ye�a:%�Ʋk���$�mMe��u���Ũ{�|(�����xŬ�]�b(Ŧ]�Y�	F�	7��#�P��Ԭ*��l�vSS����s'?�&��>��Bs���1����r�;�X��{�b�>�J�pr��r%g/~�ڬeE����>5�mb��T;��Z�E�}��CC8�ٴK�/!�����9$	�J�x��bg�5lo�>Ծ?b����~�͖5��+��Q[��Vi���q�:h�ȉ%}�T���kk�Bo�_o	�ΰ|�4��8A�_ �W�����{�?Q���܌Q���A���N�C)b�$�ո��p�_Q��ƞ��[��x��ڳ?+nx���f|�q�_?��Z��v�rܥC����j*b����v���m�9f<��.�;0�xǨ_|~!N������+�ŏpN����X�k|�WJ?�h뭏U�O��|���d�|�%JF�k�3�n�/�ޤr�N�6��v�s y�-�
&`Ż�s\K�C�+ͺՃ̝�[�!��d{�zS�V�¿H��\}tF{�˘Y���Z�!U�_��{ʵ^�r|�ԏdNS���ٛM���߅�d��e��j�/�?%�D0I렽|�Y�t�%Tr���}��j��OE��be��Q��;��A�&s�@�z#�^0��Q�R;O�%�N!�l���ӒV�HM��HԿ�ژh��^�K<��.���+�[e�W;-�a:�d
`��0.:O�E���&~��]�U�,;���.|�.;xxe�-Y��/v7���M�9���q��Q�D`�,� W�ul�e� v���O��3Ƒ��|8���e�Җ7�:v��|n�t��SsPw}��|-��/_e��~��|�����sܜtg��4��M���6h���WB�?2x�}�Vu�Ӌ<�׽C���� _	�<�O_��[!�4���yK4 ڸ�z�:Z�e	�H0��~[XK�9ZS(�	�4�F�U�%K&jڴf��`&�ɷ�۔��$<S;s��4��Q� (��Ds�0�o�l?2Q��j�U����tK�5\������=\�m(�[��ه�\�����tB?Kyg�
F�~��~�s����"�kYT���U��՞Rs+�;5�6�*���F��!{i�� ��Y�S�N�����������E	�Xp�����-?���\!}b� ����DŪ�=׵W�����尤�����׮�G7�4ʖ7�!'���yE� ,�}��&�܅k�?��J����4:��܏�e /���U�<�12!T�	�6���*t;�#��].6k����Y���fw�M���b�z�f�[������6;W�,��t��ޜR�,7�&�!Ƈi1�Ȉ�O��|*�рio*1� ��U��W�w���+Y����C�W�x�g�T�:���[R>��SU=�Ъ�=zR�8��ɃhK�a,蔱�*Χ9�[;���c�ø�_`�l��Fn=�;��+D�M�]x���@�3���0-G� ��4�P܂�e̷��L�I�A�N[	!l��؛�!���"q�OB��a<A-�_�8���p��ˁ>e"�q�N�MX1ᔜwy��iq����	5��	�,�$_�2���1	eܑ����ex�����W����F!�Yw�5y���Te�L3�k�>E�����~���m\6�q"�х�`���㤓�.���U!]Y�ɫ����w�8lm-֝G�lDƃ�0;��f6��O�����3���T笽ETW~��
˞��C77v�1"� ߗ��A�"���S݃u$P�5��3b�����Q�g+��������@��Y�2�d��#�:S,-�HnA�
F!,޻��R+%�f�~�;ڣ���]��KK}�K��~�U!,�B���r,�Z��hr�7�V#�u��6he��F��[Ea�{�U�����`耜GِVٚ��hu�Ɗy"��H��-��}�X���%��+R?�wd2˩N�����s/���U���Xw�q�Rlh��4��k��a�E
�����ZE�MȜ쨸,�ܟ�b��׳6J�0���2�NAL�!���`t��!�)I����b�Vm%�} Q�'�-�n�Rp���][��Cl	ɳ�
��:>S7�����`�5t�I�G��{�n�(�uH�]��wPr�̡�bB%���\�Pm�"O2��OR)�i��,��"`Kk�&�4	S��K�X���n|�>c�����Di�T�ժ�Ż���	cXѮ���h�1'$�������\���m��^����?:�+�#j毡�qeQ��L+5<Q8 !��p�_�*5a_�E���x�������-3��p�f���j���aBxk��ëi̬�s ,+C��21co�������Yh_�������t���]�`�����f����/�3�z�ĩ<�%X�)��F ��قh�i���PՕ�S�P+ ����֮2/��W��M��P�>S[�iĝ̣��=F?6^zd�-�8Z�8T�W�vN:�"of\���phl�:�a���}91M���"?�73o]�mT��_��o�І��c�(����%s�32�����!`�7+�� �I�M���?��t��؊~��b꽔��Q�F�~�eTH�ж���S������)
��)�ojJ����[Dr��w��	�k�m��!�3A�Di�O��.��WDd���+�B��2�
Z�C	[l�eP�VORk�l=���6q�۸S�X'QMBL]������^��7#S����r~Y��!j\eq*vY,��GOoy�}�V�7��5v���E1p�� U���+�3�Ϳ@5�;L�}�z�'b��+���_{�`���>	D�ɞl\��+W���"���C+nT�_�>����Wr�4AAF�$�W4G�ej���{��(:�K�)��^>��}���j��о�1j?7����I��ۉ��E�� Gkן�H��X�m}/8(�5�0�B�߂�B��Ԫ�R#�>(-U��&�7���X���K��_4��-t<s�iB��\o�À�Z"�2�I�K�%���J��U�����ky ��=��Gҕ�ԝk=�|�ӛ���`����"���eJC�t�%X���\ӯ�Un�(��n�.u{�ઐ�wS.f���;@�9��~n:����UR���d��f�M0Z��^?�FX��j�x���d>c�Kw5��Y�tEk?~�j�g�+aǧF��ju��k�W��p �pL9�ŉ3�Ƃ�f�MW߻Fa�'��T�/χ\/����.6d��K����C���������'�p�=�'5u���sB�"*�Zx"t��l���$>�xzA�o�'A�s=�G/�;P���eɰC�B,%�0��8�+��LQԊ�98l��\�l���5+ ��i����e�+�	�7�x��IE�f�
6�!ċ弹Z���P�����M�78�=���h=g�����7�-��~���	bBm����iܱ�jE��>ׄ��i+cMf]WH�tG-e��W^1�fnze\ �?vp��iO����**��"(� ��@n�;hWV�Z�յRx�f��/,���7�aּ��ok�_��2�Q�+Z��jYŰ �h#F�(���0���C�`g"2��ސ���XV�ro��Y���M�,$���{Q�{N&�7���N������'e|�@CP9�T`����%��5�>j����Rw޹��5�c��Ts��Ί��͌'�_M�H �#�Vɠ4'�j�z����2N��S] �t`��I$,�؊AI����_�xVGw�������	N�;y�<�yU-�D�zy�#����=?`0 }�t���?����)2|J��:%1̪���V�Ӟ@�e��WC�������3W=y��	<�ɯ&�JϜS���S���ha^���_�D���ل����45���Di�Q����/2�}+6a�0�f����~��6l�H8#�wε9�+�T���~�y�h�s�a�ܰ9u��:�����rG	3JM�]ռ[,�D+r�}+v5_���>����q���3�Z:):+���~�K��\ȃ?��_�Q;O��'�:�F�]�J�#���m�7@x�"ET\a�P�,*�L�-}������]81�<V�����d��a0[6K���?���m�n�>}�0���N�I�-�I��Mo~�O��S�l�2~O�Mtt��|aH���d���n��������>��O_�d��Jm	s6.�����M�z3��5�d1����1E=?_�V=Z�g��4�e/��1�� &����Z�U��Dz>����@�����|�3MӬug�OƬ_��� `����h�PB�s+.�Q�R;��?`4_�@�')	����S[ȵ��ja$ G���5����YH�	r`�۩��#���ŗ<$��#b�{���B|e@��i��u�U]�j�R�C����}ejp@��j��i�p?t�q'FXF�~��y��8(C���v�{���b��7�z��ۄ/EB\��.��[�c�򀜫%Yy��	��ԝ�x�2�)%�S^�@��̎QN��a�e��r�aݭ^J�͇���<�s��^=�t���A3�'#m��4:xg�u��q�.}��d|TY+�r�Q�6Ƅ{.5lg�I��
���_q��m]��]ؕ1���¶&�(�zm�%n�h��ؗ>r��p��l5�6�Z�B��k�	����2]�#�ݨ�*����*�����ŉ	�'ԢY�������8���z�R7�Z����iJ�	�Ma[y�g�����ך�����e�ԢvŨ������dsZ飝~��Ί�*�e(��o{�.��6f6N���[�!A�z��Z��M��1?dm��S�6�O�~��Qt��ZO�R.GBU9<�c	�nC�m�*�睟�~ӳ�/�=l�um5|�}��<E`�n^�T��a�y*0cUg ��죲��r+͸�,��Hɖ�l� �������P�=;�l���Mxo�Yٓ��egN3����O��>�g���ء��ﺰݳQ�OK��$y��(CE�nmR=#]2#^��[!݂�o��<����JȈ�LzV��5�c��s�� z�k��m�x~=/��x�-8��e�4��v�a��k>���|�a��*�"�����J*�O ��(�R/@\������������!����D1d�O+%���䶯ψt)ٖY��I�u�vvڔ��q�mW~�lLA����P�\�
�O���i�p�X��t���P����yD���i$]�g͔7�2;H��y8r�S�v��@	M���G?��Y�Z����8̗m�4������Q�Q�����"�v9���F�M^�;c����
 �	�qZ�'rr߰Y�9����M#Ja�~+}��Fm��ܿ�m[z>�zi�*���&;>HS�e��L�U`)L�k����L�ߚ:��3]7c�G�[�q%���ʨ^F��<s�8}8g,/;�� A;�z�X�'����#[4��B�C����'����aT�=:��k�#j�a��׭�����7�_KtuX�Ϡ���T7���W�q�� ����-V,����(	�*�F��t���w�f�� 8_Z� 7��4�-�x�ַ��}��f{�1���+�0n��f�q�^��)��B]���J#���A/�v��O�Ӊ�n;�	�IYkO��&<�f�q�I�p��y���s��T8T����%]����;�����UD�>�%����$���n�C�SP�NA��A�;�k���~o��?�r�yf��9����h8�`���U�Fg:��U�)'�_?���B��E��$�����nQ�Č�V��Et:�fa��{j��k�2���u��S@v~|�9���vZz��9<s̪I�������u%󃥐��CʩԎ�=&�@�[󠊂7�O}�� ��
�\z���hU�̝a�Tb1�)��}�4�Zl��$��Ky!��vq/,��Y>Hv�9�)ZπzX�C���B�M��u���c�@(�M�)���s-9m��q�V�H~׾�7��(��k`���Ic͇���`�T���kM�beP�@M�yH�V�&~.�����q(P0V��%*�1=';�y�p��%�d�U5�	�C?�W�3��6��7�.��؜�F��l�QR�T�Jag;Zӆ������|_SkǅS���JBV%�K����"WL{���������3%��|��.�v��,֤���Rg��S��	�yVc��P��Ƨ�WRe%O���Ԫ�7B��Q������5Y�����2ʞ�^a]�n_)%a����ɤv��I��5����m��j�YwS�@���n#�l���Â���`�6Jq�~cѨ��ȝo����,J��a`��'[[ķs����)���Fl�j2C�mתו���L���J<g&���g(�X���Ϯ��^�]۝�5��^`���$7���,f呔w�F��0KvE���X����ͦ� �ke4��n��'�{����ۄ���ӎ�-dᖸ5c�:��|�,���w���k����U��m?��V��K��(��zx��?A{vt�3�%}Ѥ�3W\�l�����M9���ٝFX䨗����2>�L}	���u�c���c���T�FO�����[+�&\ � ��>@{�"���y$�	���)Ž�����G9�1x�=.޵�9���	<�vo�U}��9/S�����i�!�yHYM糾Ox5�A
A��E����x#�oM�Eb���uL�wj���笠4^?�Q���eT|�A�G���:�ޫҒH.��~4̏k?%m���u�U:�u`���H뫣3��ͯ�Z�Oo?�>_T�y?#taT�e�D��od79@�AU�v���\}�EK%�n&ڎ��K�2��;vm��g���A�n�#���A4^\Dhx�R��Ւ���g��Km��Q�΄�^��y�x���V����$j�\��.�ћ��G��2_4UVd�54w+>��W�Nv�_����<6��������7d�ٝ ����b5���\J��z��Po�9F.���V�P"s���x|㩟���Քg�ri��)�B�^O�g�_����#y��ۖoЕ)�h��}�J�)c�Db��b���t�hU/��OnfsC#�ZjZ��;��̦.��>/�U�D��8�F��U" j�3Y7m�1o^=J��ׯ�xs�L�D���"�!3|˷z�NjѺ?C�p���ZZ;�~�[��"r<���*|+#Nx˄�L�O��u����LPѢ���v|��?{2Df���2- m�G�\DQ��ok`ա�ʯ�Dc�Z|ь�^#�m>u|���Gb��q�_��|$ꩅ>XK{�I��㵣�$�/6�$ۖ��0�K=I��q3Z�g��2A��J����Sg�|�w��IT�A䈐� ��w�]����c��űO�?`�z`64��sVE)>Cʭb���a�ԟG�>�|�h���5�N�vLu�o��i�~yR��bDN^l^vmD��F}@�+�Z�x���I�@ԙ��� ���a�zb��Py|����Z�x@���[�wO����H8�e�^b]��b(��5"�R��]ux|{v�&?J�������^G���_Ӏ�F�q����vP�r|ٴ哀l	D��6��
0��b9��3ͱo�b��P��04^�h����P�����_i�"
��aH�:���~�)�4� �d�C�t8R��<�f�#�q@J�0�{�����
,��Uj�����Xph~
�^2��S��2�o)�ѩ�{2�!��D������>eYXğ�>�D�>,h�̂~A��V#dq�Mh�hK@B�w���v摒|:_��5CE��>�m;�M#�3K�U��AܞR@����B?�����+�(��
��笊��4V��G����DɄO�����OʯVˁ�LH������kZ�עmِ{q|V�<�R�%�%Ҷ@[�+�����M�H�(;���wGZN?�D�l��
�z��$�7czEyw:wl+�/�������m��#�_�g�a��9��]���@ꨌ?̭�"	q��
:j�h-C�DE��� u|�Z(,7|X����T��&�����������y�i6��ޖ�]��|WY�,�^�N�
�s)��`��xT�(�"��k��L��R`m�;M}٩����G%c+K���Tz����,��X������ǎ�i���]gMTYt�5��Q6�J�/�Z�t{ʰ��7��e�j����E�P��y�S-�ܧ�Ʀ�����Bi����
�׍6���V�m� �:�[H�d�1��6�D}ѐ��gA�O�ړ�Z�JF�?@��	�E&��4y�9R0�(��&�M#^fgX�5��!s
\�?�L�����ߍ1g)H���3�L��F����R�m�_LM��#\ O)�ڄ����mWVp+`�ߐvn�*UO��L��gD�X$!�õ�G�j��c�i��9]4O7i8�/��5M�]� &�Y����*��z�'��W�l^���I{�0�E�t���2%Ҷ{�b�f��G���r�
��\e�B�%~���Z�ax�Rg���&u`�|���%���~��x4H;�g���vB�C�UT�ج,�._#z>�*�m�/0=���QY��&#n�F5���`��}$t�s���7��F��e�b�TקB8(��Fg��@�(�)8�4-��
%;����ˌ�?7]H��@+���,���Cpwv�����m�В7.*�y��q�6��ؔ�藉�J�p��M�V�)x�n`�F�IZ'�]�?/�	�V1ԝC�� ݧ�F|�B���F����[A�l47�˽&���w�Sc�[��Smx���<��\�uJ��9���t�y�2����#�[wP)A����N��)���"���&.��#��iz���`�dv��%�'�ئ$��jC�cQ�f����l�m��(0�n�/7GS�K�d޵���0�F8EbP�����-�	��+?I�p7�@�fO����d�5K��ð`��v�D�cK��<fVN,a��=#Q�����seN*����R5���@��L�N���'	l̋��g�V�JU��i�/[A�_��H�K�-�3ּ�Vq�!�h���C޷&�y�W��*	]������72'YG�+y6Y���*��"�W6~��7k�b�z�M7�(�a|�uv]z#����Ǚ`��f&�����`Xⴧh���R��.���ň
�s�:�.� �:��%��m5����۔�qk�ʒ(�%n��;ҷ�\�F:]�������jϠ�=*��[��A,�J��8�Ð��[���Hc_S9h'<�_�)Eӂc�02�ŏdR{�vW�a7=���� �~��!�e=T�	5��7����3�¿�����#&�|��W~�G
�ZӢ�h3��@�C�vJ]]���E�{�����y�LFM>	��y�N0��m�/�Ħ������rX�c�~	s~5�{L|u�P|P�C���z��o�D���Z�����<��2+ZK�h�0Ȟ�*��� ����g"ъ��bh�����AbYX�R�qJ�,mt�`9�f;��y���N��%!X��.cXq� ��\��'q!Ѐ�x6H*y9���#��%l�^o?�E��3�:l.�l�[�ȿ��V�*�h|y�����������[>���!���^�Nsz<����X���WK�nB�,%(}b�%~�K�!�95��.�{� ���}��prG^�e`t�6�˯�{,�r��?��q��^��,�8�t�ޑ���e�_���9�)�n�*�K�%�����+��ᐮt�ֵ�_Y����L}���8)Ǚ��FZ""���6=�m�
RK�ݍ#�̷��B`gAknZ��Ú$$5�m��Lhn�}X��`�e5����O-8�NOV�����×d�嬪��R��M��K���^�D����;Q�+̐����{��U���?�Ǒ�F6����8~'��N����q��^io�|��XG��kۆ!P�uP���n}���辺F���{��/=Y�j��(��r!3��o��ד�����<�K�9b\6�-����t�y��@FPlg�Cm%�#��OI���w$����qPh�JN:'���W����`Pi��܍3�Dj�g���{[��R�W��>�eqFɗ$R��\�5���,�z��>^�}�xSj)���ۃ�U')=6�"���RNa����#�B���4�Ugf	���H[)V^����-��n���r`�ltٲ�m��Y0nOr2C�n9���n��em-0.��V��kѼ��[Z�.� ��c��1�a�Vb��7ڗ�������KI�ks�iN�M�D�PR-���Е��Ȓ�F'PQ����"���S`��x��ZA������e繦t��d3��_�i� DHe,�Nss.�����b\�$�5�Ϯ���M�x,����29�T����y��ړ�ש����j��	�x���vg5?��{�nk�lb�EKߑ�̩�+�����,3��ZZ}��%d�פ���0&��L3��|,��ɳ��_	�}C���Shx ��'�솃����j��E(]jM6+{ٔ\uP����[,�֟��? v�-�ל�`��d�M��HUƤ�p6l :0�ْG��#�!ZhiV[�C�O�+�>�{}���zK��n7����>6�?M�U.r�Uj�/䌴�����U�b���J�F��v�C���!%8�<o$�:�E�3�9�vD�d�!X^4�_��΁J|�w&.U��Im�iz!?�\:E�&4�L,R��ǱG�0P��6sQi`���oӉ]���hHn�:S\f���a��K�v��n�d�5q�_lC>�(Xx��@T%(�����`�e&�CR˺l�6��g|�LnU��+��3v�J� �1B�o��Yn�6o+��^��0����ൊ�^ ���0��s	X�rC��;h��N��ԛ��X�Ds�8��#�pb���.���9��]I�Ȓ�u:0S�)|��O�	,/����1�E�,f����1���_m����$��t�=!��V� (�j�}KEb�I�@�P�^f4�IhӔ���gd�������|6�� ���&uH:a�~H3)B��b�v�ͨc�z��&B:��b�NkS�e�_�J�C��\�����V��"�=�a}2�q������T`��<d14�e6C=�C&�E=dG�j����}���4���Y޴�)���KjD`���Ĩ�*�;�tc4�(���;\T���НLE��'�
n��s����s#�d3 �������8�S�9|�F��'��%'@TA��x=�����10�'���6!8XF��j46�ݖ@��)մ���S��h��n86��Y �U��R�����a�����T��!���M���㇞�1�+:�P��쭱v�͋xؿP����(�����Y�0c��2�R�=W��i2�7��͗��L��:�P� |<W�w��l�9�Ζ��-��}u�93J�ߨ���>ni�����E�k�nY*8M������\D�S*�ҏ�wtdNl�r��e�BU�^�^�.�_���	|��{��o���R+�L�n}��:�5��;'_JuF��?>�Dz!�C�_���݉ף�5Kե�Uz������"�w��z��٘g��9�c�Е�h��7|'I��vs�e�����E-��/������E�J{�C���=�I|qua��i-�^1��pk��Ȏ�[TM����8��6f�~ʤ½bk��R]����ap-<�����vr9sh�*��Nm�:>�-	]#�!ȶ�)����*e�ǂ�n����F����E��ԡݸ�,ˢ��>댑��lQ��lo/���ԃ����	Ϋ���;F�'��m�.�
��f�?9��n��ꕴ*v��Gh����ޅ	dG�	��7�����K<���5����\d�e�g�փ/ّi��R<�Q2�-3P��6��8J�v�ֱz�N�A�k|�'E1Ւ�d�`׭��C4̆�ۭ��1�@�bI��;�n���C�4�s΢�s4�9��M۝Գf`N��t����i�_�o�:.�����f�2xܾ��E@kjehj��������dkO��>oFM��o��6��a~x�0��!0�[�6��{�K�����g��bF�=�n�	�l�nT���S+G"/�za����g����h�ů�>���B��O�=���(�B���G<;�(���"�y���N|Г���Hg�����w1{DS$���t-�8�Q+={ن�)Կ�tW*�)����ݡ�E¸=����}��p���
m�p�´�p&��?8j�+o��/`�ԛ��U0�|ZY�M7D9U0&=���a������k���Z΁6π�W\;*�ԉI2<��O����{�q��K"e�	G���AJ����(�@<Nf�&���'���+���]]�� ��Aٲ����KTp��<;8t��4&NZy�r���b���vY��ƺ��!b�Kv!途z��m��X��6�XP3t�=��`��v����q�j��¼�%��Pn>e��N�G8]�.��w�@U��ҍ�/e$��m�U�ފ�6j+P�n�65��74�%����}_�Dh[�ͧ���&�����E%��J-��j!^�rS�9ԙ�G+�k��5�KZ_3�6�횴�8�χ�,MV覒b$Q�4�9�Z�Vk:��=����%E�Ɓ%g�Mϖ�;��A{�4�����VY�ں�on�l�/��p|z����7��ٯ�6BV_v�c�	�Mc��W�"y}ţq��{�9�[�`�k��%R\!�Bw�A���W(����j��z*|]09Ф`��f>��ՁF	���n����y�=���t�W1�њqB��b'JHJP<3{�H@��^�)X1,��WU�߄>�u&1L�?���;R��ɨ8� ���qH�C����j ���=�M�=�(�5���*ͥ `nS|3��9�5B��0�`z�<���ON�f���@�y.���E�X	�U$�����&{=U������A#M������P��Iͩ:��Wa�6n�(������ht����4:�G3��UX�F"Z w��}4�~y#v3�k�����2��L������#����ԁV�+:���]d���k�L3^츚6i�j+�۴9J������n�I�>�%�.(6�1,M$���"1_j0�AiO�J���ґ�`�[���d#VLC�ݶ�cZ%������w�ƭ�fA�eW�As������[�2B���c�]��Z�6Z�Ғ�hJ�p[$S �p�BF𩸉.t��O1���*����=���4"y;�C�!)IfE�[_U6�)f�����[��F]v�����-U8�mp�ƼS�������~`�l����*-鳹.r��s��,`��$g{��Cj�NU8�>H����7� m�`!�i�*2'o#M�C=Ιg����Ǆ�3�ϗ��:n1=�|����a �~�v�����,X!/\ҥ��� ��[q�娽.�0EW�;G[-i�+8�-�kxQ}sJy@/	$!��ZYџS��nY}�!�U��d�w�Rlఋc���n���G$Z���{uoƹ������2S�J�E�g������D�MU��#��B�""����I ��c]�H�Rw�>��K6�Hd��
IRHi�b���i��藈ic_�Z������!�|3m��@G�1�D��05K;|�SO1��Ͽ?JF0"�����Wӱ}��'�a6ݐ`�T'��AiRnX)����B�L�B\�J�6���8�Rc�x�ˣ���+J��1'�̶t�(9�����<�}W:�t�,�Gbv��Ri�	V�x̵���`��E$����=Cd|	dS����B�w.�i�3����Ki"Eψ
5�¤R��<&����5��N1�����f���K�m[z����ry	�Y�ZsIdS��PxM��i^��|��]h1v��K��,v�א|t]	�3��|2��\2��DG1W�������_[��z��BB|j��3��]�� D1L�|Ɇf�q�W�h��a��E��2���D��ӈ$�6,��>C� ���a�|<�Bt�����4	&���Z'��.�zG;���V�pǶ��>��`M�������� ��1�9�����Ӈ��A�`��Y.+��х�t�2sb��Kn-(�w�|-N�����s-0�*R!�'f�"<�G#��D�-�]�&��	�!�$�a����k�j H�Cݵ��qY}�ƈp�w{����xI��ψ�>�یt��+8WTZ���^����H��]�����$����Za��GWWPȤ�2�����%=27{Qy�%�"�`�T�s�N�ϭ��٢k3�����I\KvG>��eպ�d�Q�^��D/�$��^�o�궋��*�^��wա���>[NC���e�����=�l.�K]5��T66�ݦ��e��ҽ~=D��&�M��Sb�����oę��y(�G>�*��<u��ӣƅ�E�Sˍ L�4�����Kh�o�������I$B1��וj\�>��Ǎ�!y�~X�6�m��~�xA^vZ��?`)�7�UY�H�-�:J�hg	뗄�"L�h�<8M-��P��;oٮ3)3�J���[��݀x,&����h���"tک��N���'�7a�;�p>�I6�x��Ƀ�VJ[5L�M���٢V.���}�\�cX����
$���}
@�=��am�/	���©Ce��%�J���F;�ǳČ�v���ܛJtř���Ȭ-!<y�|_-D�~���xA�4��h�n�:o�"�A+U�2_��>������忁�t������X��(gq�@�=n!���D�^�N��fIK����D�2�'sw�Y�t�U��5L�?x2�z�ɝ� 3\���[�����i#���=���0h���q��ߥ����O`B4H�8��_Y�������\݅NV��M��ػ:�A��R�`!92��ݠ���Mp�i�k���m��x-X^^~�g�;�'�;5��"i��9c�.�3���/��A?2�֙�ԒڄDS@����mQ�m�/�9t�J^Se��-|�?��_Ǉ*�{���0�v� Qtl8�.�ܡӼ�jF�5��5{�ܝ&f[֝�ҙm��K� ��~�h>�k9�	�XImo�s��w�^��5H���t���k^����D�6�wJ��� ���0F�mqX����!�\�8?;|D�����kL�y�d3�UYs[�YVy��v��5��W�F�4A;b����\W�ak���^H�pj :�12p�b�١�S�����d�jG�Ys��ϷG(��ڍL:�oo]��Y��c;�w�WP%�)�?K{�T}��������學0z=I�6��o�P��l+.��ɀdh�{���2�����=%A�"��%�
0������j&����r�ҩ�(���?�����n�J0�q��V-���-6Nӆ��^9��`�o���m�ZKM����I�a߭4�ϲ�+�f0d$�	W��SP�c�5:�c�0f$���,�k��Z�V\�y��읆p����W�����z��0cSB�k����xBB �����'����(�GMA~b ��g_�&[��8�������H���^TD��y�tS�Q�s,\�1�6�nQ�kg?f�qOѱ���-��F��
iR�Yg�"��%d��m��@t\�v�lnh {�y)+���E,���Z��;�~�w��M(գ�i��鲚��E�*鍂$�Π6��9����s����v屷r��1x�R�(�R���nZH
�^Z!x� �Z����W�('�/��r)[��n�ۄ,)����^y�j76��x�^}}_�_B�E��>}@�ب�f|,�	���_�ϰ�ۅG�#�6$�(�Ev�������Y�E�~�j�s�l��][Nv�n��G�/߫E\]�)y��~Q��d^智m�S[�U�o���������pW�WȺv��-v3� �XW��rzKdE�'��c-�HtH5�Hw.�/r� ���T�!n@7��ް�hs2)@��K��(��Pf����O��+4�;Qo
�(�G-�������nӚ��m�U~�>0*-¿������D�ym��ph[����M��󦹵 ��Lv�;8��p���۽������!o���f���ҫ���c\Z�A����h��
��_R*\;w�����;�/N�B�x��ri�4(O��^�W�g�-z�3�fH�X$�Eٌ��yg79s��ӱm�UM�Oc�6�Ɨw�,�]1bh`WR+�Ƙ��c�]��ο������d9��Qh�34��Ȟ�>���bC�=B�+�-�f(n�D��V���+m(3>� s�:��=�������:x }Ñ�I�}�W��/�/���_�����6V�ur�twJl��+�!bN`��M�c9m�dI[���}��_mQ���%Lǋ���~�_�4�:=�������Oo��p��V�+T`��S4��n4Þ��x��^9>Ǽ|4�*(�#\Gw���q^�"��9���M�8��6�����؉Ij !��ʌ���D�a]���!	�ر�J`0�ʖ�fˮn~C�P�j����Z���y��qA[��1}s�C�/?ǁ@��Ĩ|I�y҅_\7?a�CX��#S��m(��'
��y��~�?��8�h׋��0=H�f��@����1����Ex�J�>p��'v�n6���T�+��)wA톗�����������h��99�B�ԬW~/�:�e�G��i6Ue�<��U�6���'ڂ�j!��! "�W�D.�� b<��RY ���Elŗϛ�֟�T7,��LB��eN���r(��x_���Z�~-��%��Zw#�K�,�Zl$�i@ip|�e2��_��	��+���J뫉�*��K�Z���}:�E%Ǡ���=�9o��A���zۼ8F��o��%���N2�)�7˒�F��*�����|KAj�uV��`��n��!�O'|ٿ�^��V�n��+]f�n�n�~X����N^]� �}i$Pԫ
����B�6��PŴBzd���`�:�[H�/?� �poLP��B���E�m��|�ϼRT9E~�_�	��o<a�B��D�ԛ3��v)����ڵ��9nN�&�4�o�:��s���.�
H'KQ�-�y�?CNX�n�=Q�c.ȚK�8˴�y���*8b������j�ҷou3p���vN��
��6߾h�:�5��h�D�1�d6�C���$l׺)1ŸF��%�h0.>�
{��L6	���\��hr��B����13�ߢ�AI<�ұ����ϰ��2K������&��y��g|����ǥ�`�BFP?�C�u��AL"S7lp��B��m���mcJa{��ry?�)>��A�7Bf�M�����ODӮ��w�ڨ���B���7`ݘ4:I�l8#̐���5k���y�샅������"��$�PO�$� ����~Y��f!���cp�4ԋ{�*�������F�J�0dp#�pF�1/:�:�J-�z��%n�|�ի�-HXTa�K��g�_�]�x��e4�S0���5�����ˠW��:�����)1���_�]O��2	0Z�c!�;�Qq��)���9�l8Rk��|�-��>{�9깎4�^T�v֙�\�	����wmu>�y��c"��m������t�/h�{}]�Qx���)��G����H�@zU�n�u^����u(���[]Z����ɎǙ$d�Т��k�<��W)�����ܹ٣&2J���j������>�����7�:T�Js�C��C���5S�7��x@�U���R���7���^A�N��|������+'H[��S>$�'����s֋�d���-�1+�_P��~vk��&���soz���2Ρ����!sm�A���[�����w�����w��A���t�af-�E�O�l�}��Z�F�����M[��8m��J�"�܁��:�r؉j�'^��t-��R���`��'L�lk�:]��:�����4 ɩ$E�/��dZa�3/����'>�$��C�d_D�I���)>j���d�A���X�)rV�J�a�6���:I�����8��+�-X�r�9�I�qz�������a6�tDh�J#ab*2���2/�ٺ��5�nH��)%0��d�ĩ#�7`��AsT�q�b�G��u��3�3��ĤΔ��)aG$;9�5)����_�/�V�d�K�;����u�؏yPh*�:��:xl��ok�y�l^`UT-�Hԫ$��Sy}�n�)����I�K�Rn��+G8'�Z锆�	�	���[fS�墾c$XBz�l�,�`���O)�Kd8u.G� �0I��U���@�Xx����01�b=�̆��2E�ѳ�{?}��΁�7ϧ��;Շr �WԡU8Iyo�5�

��(&�ș�U��Z�:=����2�u��O�;�v�&�.';I�6��]m�]�M��]!X�ؕ�"G�]̳ߤe�w-m"�蓗�c��ؿ�Jvo�[ﱏ�Ǩ�mB�F���!
������}o��J�,*�*g)�ʹ�_�f>�B���N����(����ؾ��_2����V��ha���i[��$��or{�x� �Ⱡ���a��hA-��m����R-
�����<N�˘�\�`K����Q<��Y�H2 �9�0OL�gPxh����K��KO��J�9��7���[��9�SP*��=#��Q>�������Iy��wo�,pw��aܼ��=��a`*zZ;�����N\��9GN�>��8f��;�^C2ߞ��_L'��G]7w�{��r/M�[���R�$�.i� UP�lX������7t�1�Ѭ�v�u�]#aRl�]1��:L0�ա��V7���#(wp6�bH�J���][!kI ���%�ED�H��݈�y��f֥칆V���w��ľe�r�Y#wa'	d��en-�s���)oq��K�J�Xa�#��L�����81���+�Yʣ�k�$���N1�� XS�s\�~�a���YfkKPa/��.���1�����H�[���م�����x��;��P�hpg��#'(�5���?ڽLp���X�_"�&����0s�D�������H�k�"U��`���΢ѩ��c�8��_�a��x�Ҏ�8��¾��������.5��(�eac�q"��X�`猿O���*o(�#��i&���Z�܉��/������ \�:��<7Ԕ��.Tz[�0�R� �YG�b�G�V�DT��'��Z2�(̕� ���{���5�`<��͑�H�A�7t�n���D�I������
��s'{���H�S$�?w�X+g+1�	�,����V�b�x�@�vg���ˊtC�W��������?	L��8��4_7��8��)M���AS���M@���<.�e-��^3�V�����;���#�}�X^�Y�����Rb�{w�6O����g�{ޮsb8Z	�xg�/(�)Y��!9Gk�����#~��`yj{�?�bg�)ha!WR��e��2��9��H�Y�.B�h�!�����͔(������`�����6�> _�%��v�k���&�����DP��߬�q�w����";�����)	�����~])����u�↿a���j���AO��Mڿ�H|=�5zoUe���oD��q� if��k,�*�3�H�N�������LJX&�������-0�^M�l����JK�^]�x����2�C��H(�]����ᵛ΢N!6�?0�u�;@o����O�XBo=�e�K����[C`�,���N ��z����da�>��QP�>���J��A����HBk����?�03/ЏD����8�W��ED�#���ĤK{��-�|,���?������J�-��%���?�o��uGӧ��Ȩ�ǯ��1�����ˆ}8B�,���ӕм�c�it�J{E����7Y/��nր\�?�SlHf�H��q��LOdy0����'�mP�a1~	&J�y�?����̜�}��be,��j=-ݼ��"��I�#�����0�. ��Uʐ�K��Mz��:9Zb�N��8'Y�܁/R��G��+?a�D�����K���{�*e�`�<!�&M����iL=U=�*��ՂGr�q[�]�G(D��f;���4t����*e�*��;q揁D%	��C��uYv���V�l���Kd�����z6��k�h<�α���qE)�Z_��q徙h+$ڊ�u��
��]<�� ;!��"1� �����6��P��ɞ�/H}8�w�2��F�y���fvܧ[�9f.��(NT�|�j��~F!�B;�s���r�'�g�O(�֓��jz�����k�to5�=9t��i��vN\6I{{��6��i+���Oe�����9�ӽ�h��J�#�n��U=���&��:ty��n��.�<�{�}�b�r �MC��&�����6ZCa��{����:b�����0�T/��1�l�¦����)g�]Xē_"�J~!)��v�I���No��˯n���ΰ'������OEM�� j�ї�s(��v�����j��J��*�u|R��1ڟB']����}:���%�}���3J�u:y^�0�J}��$I�����`�!U�P�d�"�t�*�h�A�2X
	��C�\��ڡ�\�=�����Z�ҡ�q�mn9�����urňr&Yp��H�wGO���&6{�k�˔����.���5�L	��Ij�6���Gm��c�*J�o;���֛?:��}��c��ݞgs㶷�݇}!����N���3����#����������X$ϣ�����K��]�湺�ߞLѿ����|ƹ���%�b�������%I;(��
��\�u����X-��e]��%Ǹ��F�⛉o6�|�}l c^m���h�rT9�V�K���a�m���4Ց�,�oeEW�3o�gc���J27߹PW|ډ��ߣ]�;lNp�v��Hie�Fy?l-�Q��� ����	����mvչr3>�a�����2��`5�3�,U��1w}W�]+�RT�_5W'��W�����$�� ��Zh��l�v����S�|me�D:|S�)�kX܀l�h���VKƦ\�7���w�l�:6�X��Ab?�ʤ8����-��^BD�.Dv���O��J9v�"�"!4�#�jU�Dtv�V[������l
܎�J�u��|q���HW�ƅר�y��֜���q��t�9k�`�F�o�5 �$n��ر:SA�m|����\����A��ݙ�i��]$�8��(��27�R�2Zz_f���Q��f#���?T�J�,�m�f�~�f���#���%�e��J���������ČzmVxe�o�"{�R�K�^�p��fg���KGo5�33Kj֩��T'Q=�һ4Xj6Z�X�a���]�;���m�T��SD4���������o�3t���|��gQ-�`ib��Oɓ��i�w�!�=tT��ފ�K	 a�ۘ	\��Y&���SL��k�b��h��J5Th�7[�a>9H��*�t#��|�_4d_g5���%QM������φ�!UI
2W���D�(���Ю�{�3�t������3�%%^T����������t���'�jܪ^�y�W%h��>s@}[@"�{8h�'���V]d�S��mͥ����Z�#H��^��nG(u�� �}�9�`d��#ܾZ|7����\�!CG!����}��>F[
�Z�T�$�M�`�3����Coo�i������ѤT�~��y���P�k[�#/��� �Uz��]ҧ6��&j=�ߚ���Z��_7�B�Lc���U�7xo���ۨ�k��ӎ]V�i��w�n`�h
�kE��O�澬�k|+�I��YG"�|"'�F��,$��3Gh�:��-��Nr��cZv��q����M��C�Ʃ�˘�ʼ��=�]A�ǰ;�g��q�+RdF�sx�5�꒩��,+�eo�S�<O�+��<+����5�T�<z>�&Y��*q|Ғu���s��imq7��ZoQ0 h�GW@�JG� "r܏�V�è�ٵ#�\9�f
"j����s���a ��+�@�!K7Z�S8�����W2��yȄ�HP��-t����]��ܻxdgstnp�?w�u ��FM+2c���E2�]T�U�����wI/i��&L��yKip�!�&Q�{s,���9�'P�*�����������JaT��=t��?���0��}2r4��S7�}�T����k^�{\��Cry��堩l�H�З�F?��d���Ɩ� ��`Y�5��սgr>�1���^�����Zp�)�1�g��W��'����W���%��{�njl��-����0��v�Ê$�|m#U��UE�ػb継#��'��_Q0��4|eT\M�-� ��L���������w����0���ww�3��Z�יuz��K����9��8�y�O���v���כ��K�s��]����تh7$rP��N;�L�׃O��S���
��Ϫ\�96�}2�\v��MR��P\���ݷ�=�=�]���Jz��(
>y���.Q���.�'c�Wg�i�h�S�� �t=����-^�P:+{}����HYB�.�6�������DT-��o�|M<��`��o��̷VԻ�������OO'V��6��HU���&h��>׽'b��)AJ��938nY�<�b<��N���8�[+������Gx��놮��FWL���<�)&V>k(���mh��_/ f�����;����}2�C/;���au(5BAVs��m���ꍈ��~�I󞰹lb�5۳���'<w�g����m�If̉����3,������'�<k
h�uZ���0�����V��������]o债�;mC�-�`��� ���&PY�J���,�Ͻ8@��'����4�7����w�sl� ���g��:`�-����:�]i����7k�k. ^���G`�W��y]@`%���uLX� P ��	�4Ce��û�!类�H�f7Av� v1z*��WN���v�`+��y�* ��6�^f�,"�#h.��ǰ?WP����&�v�^����2�����͓c<���d�_I��������Q��bEKkv�*�/�<n�(s�l�e����wT�h�^T��������$�}���I2����zf�ksg:6dL�-X��;<ld�{��s����e���j��	��q���n��O�%����8��ܡ�䝈� S9z�8���ô��2� }���
*V˵"o�ыr�2��_º**�]2k���8�D�v]<�����F����+���{�U�V(�	�6����8A�A�r�]��n37�PG"�h�!�8��ݸ��y��� ["�?w��@Zթ�ʟ*�5���� ^z����g���C�t������)��G�$�e����Y�ev-]yK��H�͉�����&XkW��WՎ��`Dg$��^OW�H)3տq��=�.�K�qO��09	M��c\N��`0��TL$�K�T���\������&��r?���x9YM���44�biG�:ۦz���x�D��!~0�Q��Vo�7����`��l�+oӭ�R;���AH̳2=F��ШD;�hx���#��ۼnlM(r��ނ�
3���a�����Zn�����^���O��|��}L�h�Z5:�JJ? �-��d� �B�����ê���N���}���n��m{j(�8)}cGYP-�J:e2H?6v�T�W�G�&n�m��ya�V�@��Ǆ�$�S\0�ܹ
��<X�8?|�"�
n����NOZ�<��u��F�9�?#E�����O���"�K��`�)�%��e���@�#��~��I2eԤ:1�T����к��j��c5��֧�x��N�8)g�(^0 @�I.o��jғѴR�fx���u��QSu�~�5e�n�������e�*C������k+��P)/�9��K0�����P

�e�&x<q�7���a���O����G��Җ��#._ٿ�07v����� �ώ���gA����YU�ߧZ�K.��D�Xg6S�L��k��s8��|�N�D��C�~Q<o��9��^|C�G-��UʆW��m��J�Qsɱ�¥�~�m������+{8�����0s��[^g�I2W�e��<kFv�L�ڒ��5�n�^�*�.�P]���������/��<�_�{�C��;��U{n�h�?˒�dn��R	s< ����8:^�C��Y�h�7�=$���Ӂ���	�ڰ$���:�-}�jJ�c2��^Z��)�V�4�C�\g9��79�]�=��q�|��������։0��S��䩮	��J|,t����8�J:��A���aD+vvZӝ��kH���_;��ӟ%�M9
D5��嗑jQnk�퓄5�2��I�.	�Eok�,]�C�Z�v��l�����( ��<���kBA�/��91<]����[ѩʌ��+(C���N'�&��%�%x����Jxn����3jp8>�4Oے+L����ߏA6�:U�%�SKwT�ב�M�>w�,@����b[
�&<�s�!W�����Q���M����j��g�g'r�@Y$��ď���[@��8�<W��W��ȝ�1i>�V��>�Z��\{�98�,νƹ[n�yd��HS�����4����GK��R�mR���]�=�<9��a���.'|kD*�>��)D2��f=����B$#�х���Ӗؐ�L���ׯ�Pԙ/�ȩ10��6W��Z��vC�0<�UX��x6z�C��h�JYf�\��/O��z�F���F���yĈY��"��'H���H������N���C3}��@��ibn�.����*]�MX	P���~�ʉ�kj�R��z��E��A �Y:>>r�ɉh~���w�{�a����?*hO��/��8�w�`>�����z
#�ԝ�R]2je\/Si�KA0h[3��T�� �W��k�|���FG��a�����zS M�1���zJQ�+��̹"�z�%��M��0>3�\a�MY�����<���o^Ǒ^�gV/B�.h�s�=��<U��f|� y�0)�0�&��L���G32���RR«��Us������D�FL<���M�б�h�w0A-ҵ�[u�
gp�ļE��A�K�,dn2�C����Ne�j�5jG/H�T��Ԓ�r~��^� �|&�&���T��L����X-�\*��Z$q�iEMq�]q~R�N2�b���Fv$ _&�C�C�Tcy~�6�Ή�� T��� �X-�l��n�^��d��b������&�bg���GF��ݹ;t��	޾�xn��������`�_1���?"�\ؤv��dk��F��Ѧ�t���)�ł��yu�?�`̢����7k��Z�ň2"�~ʭ��j�h��z�_�]B,%�[���+6I��LK{��^vi�Z�)cvX�FP3��ֱ�=ଜ(k�l�g�:�L�h�i�ވ�	ʯ1���e�����]��4v����ᩩ%>.�!��܊
�z�����xL�o-C�.w�����~�����yR�T�݈ݏ����j�2[y��"��XU�Iܰh���ǰ��3͎�E���	��nL�g�4�+���y�6f����;���"好��)�|�~٩]0�ϸ��d�F�)6;�Y��*v�ഹ檧�c�y����}�cj{�}���(�g3�O�������+(+._�&��kfzگ��(��f�)�@-R���KLc�8��ߓ�w�6�}�LaR� �-+CEi���D���ͺj����W�Ga�5A�n`'g����"Ŋ�����V�W�Jr.R�B`H�|`*����涔ک�) �$g2��c*�?�H�kYY3��h,$�FP'N^K+2��4����z�Z�� ���Mo���f-�6\W� ��"��َ�X�Q�s]
p�3�� ۸ ���os;�np����Z��4��Y��'M��9�&Jjmz{�ʺ"R��>�'Y߬^*�����pK_.��+�fk�#S+�tlZ�̧SsվSb�2�{�ea������^��\���c}�c�@���Ӽ0,�S|, Oy~~��f��ֶ��}{{��w2薻�nNJqt�.�B�q����X+�E��%���9��y�6^)���y�D�6����Ԏ?^���k��	pƩ�s�����?��[��Nb�wRk�1��)��4ݻ;������M+�x
����_�UOu��@Ax�4߿M)M	%v�ޫ�qo%~�ݐ��s5�}�1���T�%���f�< pG�[P�ioo/���ܻ[�Ɔ����I�g����f-�t�9k�7	�n�k�^)5��F�fc;��!��u��1�Ic�//=��Sl���>Z�u�
�O�Y0-�p�=��Ɇ�#KZ� I�$m_��{��Q�cK(�m�!jwk-8���0�C��K�М�#����_5��7�a�7z��7>���8�l
،Z�Ch��M]&o�Уʶ�0��e:=rI���@mgp�i!�pE ����~��]`e�.Ƒ�EEM��r�D���*-mj6ȃ��o����,�ʡ������e>�j�e���jl������ԝ��*U6��&�)��Ө�d'���kb��Y�"p� �N���/,=)TXn����h��
ܼ*�ɝ���_i�Ͼ�f_vs ^�B1oL�C#����������4sED�<�m��N;
�p�l��ʳ%D�s/]���L�DJrIccrK����nIj���)&	^�E<$k�&a��J2,���p��]w�G�����	�D?N��m<��'cͷJ޲�<5�c�^�
a=��W��S�2/�oT�<|n	��x"J�i�n���Т�&fXG��P�}��5J=�2����h�vZ�0`"�gf�.-�a��	���}wW�~��������Q͊�+)�8����՞v7n��np�^|ķ#q����M ��%H���W� h� �9��ED�����R���W=)��>v�of �Q�w��s�umN�t��
S�r4�*#H3���Ԕ6.���J	���z�
sx���^�b��ܞ�d�Ew���]�����]]|+�$ҙP�p�NB�,��&ˣX��Ʋ���x�� c����肬��M/[����bfn.���S�<X�/�H��΃�T'�v�y���2�ۅ��c����t��#���7��w4���lx����T�ũ�28��;~��Z�E*IXU��Xy?�`��yP�����S`#�%��FK�hy��Z("ӽ�kvv��
�v�������
iX%="�|����5����z��g��/�M�K �e�#�"��Kc �B�x��S�e�gl���o�@Al�L�6{DO��]CH~£[��@���oz)J���m-�a���xT���*����T$'��d�e��4<_�F�m\V�K� �`:_<�Y��8ܘT�� �����|�r�f���i��$d�$[N�O#��7n:
���Q#�`t�s�xJ�	|��&�eX)�T�?3�dS�pk��8T�?�i�7����#�L>� 
�'�M�����Tr㲭�#�T�i�,l��Cȥ����-��]��:J�zU5��=q��/Z8�'].���ץRE�~������aꗙ!Pkrr3h�G�뿎�Lɖ(T���#�{Dj�w9����I�`�e+?x�u2s>;��F-Z�{�:��AʆStn���UUM�5N��%ieԹ�T�.�(��mGس�t?��>a2��t�1��������ɧ���	�ث0*�-�O�E��Hb���Ɖ$��eC`�]�H0w�$�Fܹ�1���ʼt��sФ������@����̜�=إ���57wn�>4rc�����o��}����w�J�1�Y���Pm���mZ�U��y�QW�ԃ���TN0�������N�� X�a�� �䪤x�q���⫹�~��1�ېu�7n�I�^�%���jW�d����dG2���M��W��zx�9�~�ajJ���B12�n)l#���dË�N(
��_�'b�T+	� s�:C�ҁ9�{�`��J��TN�Q��m�jc��Ρ2�NWε���h�����(�f�}N����Wp��⦷�"�m�km
|XÆq�M�,{.
�ɉ����`u�-��Tn���N1,%%�˚߲��H�]Ȗ��n W���v�*���K|�RӪ�y���ü`&?��-�2����䜁��i� I����'ѶKq�p�1��7a�j����I]ɪ��{����������o�ԞW��������챊��e ���=��V�{Gg�r�\t���a)/c3��_Z��4ҩ	]�|QL�v�T#�:*��W�kL��D� ���v�C`��c��ܧZQ����C(�r[������Zn�:I�+�t3�"Fׇ��a����B�L��6�F�5j�1�ŝ��@�d���ؔ�c�Mg	���s�ϑ�v_��H˒�ڌ~�
�Yq$$ڿ��^XXȶ~,�&��j98�d�m��&�hqh7Y��􍊑Og�B�1�E��5��f[􎢼!�u|:m��Un3��h�B���E���\�}�@��AѾײ��訠/p�5ŧ]۫'0@	����$��@
D���<�nfs~>�D��\���N�3��<��"	rXd��2��_a*�ws3��Ύ��ŀF,���͆&��s§I� q�OP��7 F��ݘ�;����7(�]+Jc�_Ó��u{�$���j�b�x�s�[:_��?m�UV�T�I��v�*��Q��2���<��ԇ����J
�4(�~R!�<Q�{�T�O�����b>�����;(u�v�O��f<������Z+b�3-\�:N�O"BD�c:D�ْ�;���:�G����{�=�j����=�7)7���::D���v�������Z(��:�xo 茏iY�՗T��9ǉ���T��ja�����l�TLM��V�sN(��장�������G��Ѓ�J8��l�NC�#$�V�&�N�_��Bͩ��>�ñ'�c� 9`x+M�pH3��)�m���a>��ѩV��#��c��d�}M����&��D�N��N��[���)?S�~�%��N%���i('/f�X9��3�H�\I�݄��K�\��{�[w�Ȁ�LY~gZ��o�
����!P��H�`��[���^��{\�iA���V�IM�n���Wv{H䓷��3��`��3$���i�υQ/uZ�X"'�S�(}�@��F/�L��Q��՛���8? -E�ZDx�^��>nԄ���>I�o�~�t���4�u{®x�΀9m M��5���܈̓�[�J���nnk�>{!�Õ���M��'7����ux�NW�7UF�绐���{��**�����k�b�B���jV>~�;����A*��T[���3>��#�G�B,�v����l�+",�p������x�PiGA��8l��N�߰�jW-�՞2�V�r�mz���RQ~"�AR�<�^i؏��\�Q"�,O0���%at�)�hY�9��y��p����.9�D�Zh�ځ�0��g+����Ř�u,e�<�!b﫥m�2�7�o���q]��#���1��i��b�mu�w���3�m��Ә���?��1�� )t�D�g-O<�|��2��B�'�	m��k�O���@H*�#�mW{�NB��0����Tڻ��ר=�$�}|����r����Y� ��\�������΁�\��l��5�ȼp_�2(t�J;xK\��a���#}7`��Q�%S�X��.���.i�w�H*�\����A{�zaF��d���-��T������5-��~� T�s�n�]v����%�V|���,_7+����ݣ�g�����$V�%���J4B �"v	�᝺�i���� ��ĵ�j3���^KIh���߁�|���W�S�&h#nkL�:��[����,�`��>w�>�R<�5jx)J!b`a��v�PiR�2]��r����)c^}��SE(C���_/4׉�w��M���#��[_�������¼�1�랟j��f��)
���y��T�8��e�T>�]��4O�r)��Т_Q<���"��4L�����)^b�L{-I)Chӯx2St��>EqC����	v-�g�+u����'���ot�������	r�s���+Z<i�iL|�PF�0ӵ.�i��P�y������C�B��B ��"/�Ы�3���Q���o��쩌"��Mf�?��2������I*��
�;�1�6D�[iسĪ/��J$��6\���&�ی�n��x<�R��ʭ��l��˳zװ��IY�`�5QE�kY*=<��.�V��$o0�1�x3'���g�.O'1WT��b�c�ZQZ]����|��'%4����� �jv�c�B�'�ُ*��� f]U�.|C���H�]�E5��@�[;u��Q�c4D�Â��qpTo���L�*̙���o�M�ۭ��aߟK��2���z�d�V�Q���$�9l��?���
0����,y>�G8��Ovs����e�Z��9������yv�X1���bQC� ]g����Y+V����ʃg��/s'�?w�)a[�VT�h��x�$,�t�t���?�Bf��6��l�jp�����F�k�:��M+��l��g�Y�?�Hq1�9x���6������&Ҿkh�����dP�������孍�W�,_�I��6�p�<��p�|aa��~���S�]���o��y��7��-q�(�rZ��-�>�M��!�\�� ��RJ��V�VZ�����d��?��:�$r!����T<,��5Ȭ����12�K-!HǭK��-��lݎ_}�׋8����0ִ��.�b��c��H=s�l�J��-|��<��t;�D��#_B�s�Ҥ��QrW�� �ɐ�K��ܮg�a�ىɯPת;Ͽ+����Az{Y��j�&���9K63��NC��jߌ���V�1��u
�Z<��F�rU��0�)��z�i�"O�>[�cǥ��g�C}׉�Xa�tvŅb��WF����o9��S����r`{�~�)#M'�-��8�"����^�i�YfI��7�9Kσ�AUΝ�&�ǋ`�z���(o7 R��<'�LQF�bb���+�ꋪ�����jG���)��[?p��֪�j	잴Tַ�9E[�kŇ�?����N|c/�����>���Ĕ��0���L9d�w���x]���D�գ��ȳ��WxT��n�a��}�y����M*,m�moT"t�����pu�u��u=��Ծ���-�e��oI"��o+.c{��d�|v�
�0c+�%�v�Y�jIZ��}�i�M\ߴEܱ�;r1��K�]'� ��q�c.�u����y�X�;6�f���yLR>��ഋEKo�(��G����UJ?�H�E�ſ_�q ^�f�]zŋL�)p=�C��嫻�=���!"!b����m�>��1Ҋ��]i
�X��r�c��˓�yA�jS��'�U�Z
��Y*!V��=���� ٨���.~/�k6�̰G�D�}�zR�� �:CU%�@n����&�C�f�K��HA�_��p�e.E	��6S��!���̸۝��O|w
�@��T�,ǡ}��r�&L$�<����؅g
��:�{ťsR�;�ܦ��o|�w��Ԕ����
&GS'H�-�Wڇ��&o~�8I۫��1�O
�*6�KG�,���m5�����K��as��Ջ�;J3��)�r;���Ʃ&�]R|���4J�TE ��i�'�i�M
�M��$�@�"����NO��(�m�����42	o�X�L]�i���v�{�\$�O6��lb�^��#"�y�e<�}Qx���+�Z��^|u�4|�$�{��S'�����@	��	yq�u��B�a=,�X1P�St�f�#����qy�%�_�w_�7 $x8X�x]���r$���X��j���S���UU�Hi�jA�RJ�X�U+�H��po�^L��^2=��<���WN�e�t�
κ�O�n�1V��6��G��T>(J�t���3ݰ_m��)��eΛ��8&5T��A{�ޢy�A���?�\���9�2�>�T�Y�v�0^������@���5��ܭS��ٗ�F��X�j������Ƴ����W�ݟ*�|:#���?������'�A,Q�uL�b�J<	�|zSRM#$���8�}a��qhޭER\:'�L��B���`6I���f ��I��zZ�9O�^�<���N)[���ק �C%���o�8B��$	�q���|����Y��b �f67�V�P��"��7�<�	X�@�Z(ڄ��)��#�^�W���`'��O.l���1��Q���� ��������t0�&�Zk��b s��"3����[�����̎�u'��$4�_�Qt��Ư���,u�M�9b�ؾb�DxH�t��6��1���{���2�-��DB1k)��H���r�`\��*�@�ꜫǝ�-"y����I5
d�I4X-F=Z,^��x���:�R���Ƀ��ޥg�0_Ec�;@�u2sn��Hb;z��Pʾ4_dښb7D��8	E��E&M_^��p�����-lu���Y�;��H"ؠQ1T�J3LQ6D� �Tzx�lu���U�Ev�����٣��\ӿ-�M��X�	�Z�]P��x���{�G$�y SL���w�[�_*|����~��Ao;cS�>�X��p߼�/�_���C�Zߎ��cV�Oze����n���X&`}?��ڻ''��k9�$�0W(���C�/K�h$2�t�b賃��imS�P�b�������$H9��#h�o&���)��^{��+��&����ߝ^@z��1-v�8�[U:��*Jz�Y�����ThL��Q��)��c����f��k@5�pZ� 2��T���{=䢯�s��?Ɏ���i_���HBB�`h��0E��R(>�-�phI�6�&W�siԶ|-�l:I#mfUȈ�:@�.�;�MH&���s@�x�����C�҆���Μ\��a�Y�U�Um]�I��<���X���W%�1�FC%zM�"H����s�p�Α�y�j�7�����W�ݗ�E�r�1��/l���*L�Vc����w��K���s�x鯗��L��]_�"{=������[����w��E�o[(eͅ��Ć��9�.Sq���ÜB$�:��J��p�v}�[JT�P8#�b8��M��p. �p�y��]�|�y�w����B�n҆yg�+ݓ��'�"�IGߏ��&V9H\M򹛻Mw>𫩁a����k��B�i��M'� Ҕ� f��ix������KjL;�nN�;��J~;�>����m�]�-�aX� t֏f�©�85�_���-V����������Y��bi�/�TC��Z���N)k~|�e����79A��n�]1�4���:j`�!Uw�����tv�}�b�{a�ngi+�c0����P���Z���1Ŋ�iS�7o���/�v��l����vS��*^V��ΦYv@���6�:�16!�I	���j��O_VȕWܞ�WԜ��3��I*�1� YG�%�@��蒘���N�qɞ�)s� }i\H��bF�x=�1�6"�H/*Ͳ�?����xP���p�SI=��HSo<�7�-�p!m�r1K�<n�v�$bEw<�Y�\��g	L�v^��YsfA�q�BZ�D>�:�CƩ2v25�%�^��LD=�h�g��O�c����u�m�k	�*�t�����)'O�Kmk�q�T)vQ�{FQ� ]�M��&!fI5��zS �WxxD�[����r0�ZlQ3q���j�B�w�o8$u�\�&6Z�b_�&�!I�������9S�큣Q��`>h/s�.�j���0����.���E2h_VfaH����f1m��'[�W���������,��P s�"B�_�1�J2F}���x9���M��1��9�)����@LL��m�n�H�.K�LAѣԖ�6����mC����2j��UE	�����a��!U���<1���er�������h�)euZ�=r�M3��|��N�m���E`آ�A�k�nL�Q3�_g��Q5���'��Q�2N��
Ҷ-�1�����v�����]5�P/�xq��@���:��79�"#銡"MrSզ\-ϳF>���__L��h	B�7ۃ�2ѓT3�*}��RG�%Y�4YU��C����t��~@&fUs�
D2�6�:f.;���G���=ݓ�2��`�Qo������D�������;��a�ZƁ��F�_#4_��!E������_o*q����zr6�}g����"5��"	\�|-�P`[z��ڲ	v>�%*�+�T��^STM�NF�#�K.�=mӲ�T{��3&ҳۨϗ�������f�z]n~]�j��pd\� i$��%{�!�C��%˨�Y��U�<z����Y�0d����ʒ&�z0�eq�ǿ2覨�vW� ��Ic��H|<��W.�|�%�b	��^I,0�D��d��&�{��k3#}(!�:Ց��:��A�Ƃ���ͤ�'AO�t���B�/�ұ%��+���uqjO�¢��Q7vф`�Y��"a]�RP�Gn^��"��l�+�WsY2�#M��m���``�J.Og��w_y�̷��q��i��[��M��!n�1�x]��L�����c�k?���M��A���p�#�Sd�H��Mڏ�C+�jV ��D��i�P�U��X����]u�G-����j1�r=Z_��R��}���$`3�B2��g��KjNנ/�0FKn��;�m۫�yGNfx�m �����}b��0�i��D(ڙ ��;"���ץ�=כyaG�',E�I�)�`K���z%�7I�]<���'K��/kg�?�TК��f�I�1�M$K��6�w�h7�&�.a�#�)�tX�e�쫽I!���ǜ����>�-0��Xb��J��Ч��ԉ:+?Uט����ge�C���N��g����:$7rS���e���ʹR����o�V[������ l�S�r�&��=��d�/�nu������/O;-C����S�D�˗\h��[�����QNT���Ά����$sC�DsQ4J��O���~>�[�_�S��r�rby��z|�免D~�Z+M֧�?�%��G��^1xv��A�z-�\A���2�?��{XA��lp4��2��/�#�r$⢺$|����M��N�D�������N �D�>g��� L|���������h�!LҸ��JFw3��/��(fVJ9[�����L�t4y��9և���k���G��}�iζbUg��T8%��e$.i���<�s��-�oLX6@0�,!� ׉���$�!�U�	�t�����Ӭc=Y��<n�w�D�̟��W
r�pQ���!��?1���ew̌�z��!g�j(&�m;�O��bF��scc�*�F��k����gM���9 a�B`����m�]��`$)~�A���P����-�b���l.��UF�i/IK�x�I�2I���r�[&�l%���(1��P,���4�# �h��~ޫY�Z������~B����RĹ���%X����y�R��Y�}��a�M�7cn&�gةP=ě'���_ %���8'����WO�����sk�W�M#��(K&�s���O�X��L$��0�#_D����5��A��:�����]��c�����8��& g����zAh���1��r:C6�L���F5�jx����\����̷S��	�J�	����5����r�7�~�K>j��|����$�A�W�w��[m��COT{�E��Bg�%�V�;͔�>�a-���X�1k1�K��S���d�)��]����<J��`�FV`f�pv��p���e���T�ePH�+�w��K'��l_�뉃�Z�� i�} ���I�����4I�$d��>e�ڂyi������&<`0|�H�l?�	ΏBYP�[�JЖ�o�V�Z�O�u����A��?+�i^���}���$JƱc4]�U�b����K����%�[��)W�x���l�zf.ۙ�x���X�\~PP&������AY�r~�d��	���E��v(��P�ߢ� S9!�T#�4�ЮC=��<��C�Cw����-��8ķ��JCF��ɸb��,��`ұm�ڥ���|*�����nT��_�uj0�$+���ޒէ������&����EV�-��*ڌ:tV��m �� �$�i�^̅?'�^�Ǡ��cHt�{5�S,>�9���.	S�߰��?���%�t�U:W�o]�F������Rt�� Ab���.�ԯG6�'Tn%���������D[���|�Gc�n�pvU�$��Ĳ���2��������������8��b�������^)Σ�u��.��S��	g=���U+T�(�l��=��>#��֭�%#&:�kwL����=ȳ<��M�[��:��|2�LM�h$]=M��e�2e���q���n�FCn��p�%x6+��%�?����������N��q����I
���:�qK���ɚC�u��u+f���eQ��ņ���� xz��q��|l�C4���hhU(������f�xM�k����3˲�~���VV&BRĻ����@������h��'ǕNN�n�.蠡J;v�/p�Զ�/U>۴�������n�s�j��m[�o���v�ma�7���t�t@�����	�-{�n�59��h�OC*�'���[��b5���p?^x5��Ҿ �� <D��f�7�}�!-F�AnS�^hnc�E7n�]'O�5:�a{��Ģ��C��B�yd�W)���*>�1{�֒�6"�Y5W2���7��.	v��ᬰ~��9tqr#3��o*��}�h��J����9wV�5QMŚ����r �<k9���lP�:�+㭣s(ʑ�jP��'��m�D#����n/e!\,�8on��Ӿ������vź(�BY�'��!�?nj�GI�Dُ�No.���0=m�$�����_C��)��9��ߢ�0:fX��ع�1���=|��B���0^=�9��ﺡ W\`]��d�R�_�׹��.2��vB���	�
v�8)��P�".l�rߪAH�v�M�a����~\LB�
f�!�le50����q�g�A�+�gv���<������ܽ^�tÁ&�}E/�f6��6�q���,D�l~��֫��j�K���~l��n������w�����wPON����7$��H�"�Q J�|��U��L\[o���1/�/%�Y���#%W�4E&��r� r�C,����wq�`�_-����{�HٻV��zI�K'��\�OO���ߎ�%|ܬ���y�;�64"����U�u���d��DJp��($i�Ϣ����6S窧P�;E=
����>��������O�"
���>AA��]��436����?��2V��G�+x��v�~��WV�d�oV�|�9李Rkӵb�p�Ϛ��6������ᄘ��8۸'q�=����p���Cx8(e9)�ѩ1s��~��v�U�I��7��1��m�.�����`�\?��-��y(�+�7��Ѷߌ���cˁv��!���Taˉv����y�s&��b�	���
ɛ���w�#������bA��ۭ)��r�٧��{g�i�eS��_����|���G~=�}��iv�v2�>��x�1��Uy��o� -��nP,����0��8��X�W��S���z��,'�MG��=�����߾:o�o��?'Z=�-��,�1��y���mn�\�-WK�����<�Ǌ?x��޿O�M�B�b-��L�X#ԏ�~��dB������'���V��j�r$

��e6`#��t�V���ԾlW�]��I%�d_N|&g�Z�=t����l��ԉ��hp {t,}���(3zXw9��Q�Ϋ���>L�r�F�ɵ
�ß�RB�hr��Uto����3j�����AI���xVXPa�Ngwe���?��~/}��Ұ���g�!~`7a�D�|ᰩ?Uހ�bȞ�?�:��G*Fj"Ӫ�bw���,^�P����j�u&�v�)�@���#���ٽ�eI$�	��/|�.�z�9�h-��5��3rL�֔���g#������\����8:'܅,ө
���~.A�
��h��b�k�9����U{�tvo,��j�ؚrq5ǩI��;v�aDؗ^��Qw���z�����|�O��y�:LS�"7�)'�ԵԨ^>���B��წ{�נA����kK+���ީl*�[�Z2Mҽ�=��ӭɫ��Rh�d\�S>z��S�ff|���1d���V	y��rJ�>�����x�s_�Ʃ�����qz�m+�l�O��¿.��ON���4�K��b�v�ˑ�n���K�R�B�?S���������PX7������n3��sW�`]�dX����ӱ`h�R<j�`�O�����L���à��c.��y�q�g���&���H`c�}?X��%�_8J�o�;�0�@!�!��Z:��������I� �3�a>��+�O��W���+4��89wG�I�)*5�N�$]���� ���?�|S8cރ����8d/��j��9c	�yV/x(������^�`)���d6�bz�E�o�r�j�2���_��Q:k%\�����)ե��3�	��lv�~�A5�%���nH��v�V�����"mǵ&�&7�޹}j���e=LO0��͜��a\���/�p�LI��f^i�!�ഝ�R�pJ��
A�#�ֳv�n^��o4������y���=��.��"LM�G��G���>������H�:���i;}y��q���v��;�g�4�f�)���r�T��,�^��6˫$|\נ��l�q�#��ئWcP9���O��V3��z���Ǟ
m��wJ�,#��^2dHR!���0Y���&\�p�F�l��VW1�X%���4��=}���������3�s�������6�L$��M�{	7��<g��Y��c}���Z*�*����N����#-e�����n�Ǖ���Q����Z.Ps�\l@����'Xs����Z℟l.��� Q<���L��64�8H�q�n��~6��rS����Q1(���P��I�鯌f9R���m�yU���'ʒ�^�:��<��}�p��*�@��UF���_ ��O����|�:$�`����Θ�� �(\�Uw�9���AeMv��j�g~��)�
#v�S`)&�x�-`^�j�՞�h�,�d��Ԥ#�U2��Z7v}Qǅ>E��̷؞�X�V���i���WrH
^�#]"��8x@��������}2"L'�+m�%͊*�^d�H���r5ù�6�骜��5H�¿..e��7���hq�c�\����.�w�t��(2�k^Ť�/d;���DN�֊��"�hn��v?��׶�|�:m��:�f��9t��M�~(ƃ#��'��1!�b��7�E�l]��x������^��	�/z�i��,t���!c��y
|�'9��!���z{" m[Kc�{47�ɸ�I��U��~�B^�Y����I�~�\�)v�@]e�J�ꮃT<9U��X7B���MQ�ڙ9�N21p���/��7@p���4�u��JN�h��1|�~�ԪX�DO��x�N�A�T���l�-s~-�5�sH��T��\TќY${q��9E���E����#4�b)�P��N]KnIٮ��X�^�&��@k����g��ly�q��KYaHN}�}*$�Q�n����G�n�\u�`f)�K?�\�?:7��w�=����G3��KH�~�O�*�S�;��r���c@x��)J�jl���Jߡ������Н.Д��X�:�~�r`Zp��f�/��$D+��������CZ\��w��9Fr���ԽKش�?���KA��jq�RuFn��
-��]yn����'-3 i$����X�-$����e,,�Td��^�Ὧ�բg�2�K��`;�Zb�9��S����������YB�������$Q79wi[�^$��5��4�\�1+*���?b?��)E,ߥ%�S(��_bV��|�B[6�h�\���;�@;�ތSk/(Z���� Pݳc	$�n�T��+��A���N�s�MmKk��j,���F���A3�V悂����y]�7����g늦��Lv�ߚ��	��̍ԩ�@��\C����6x^.�m���b]:b-;|��Wb֪#Az��0P4����֫�vUp%6�y��Ҫo�d��Z����Ό񠳕A{���{ğmMֲًp�> *fs���]�?��ȓXC{=ҍO���ډ5�W/�\�-.���B�wڻt�����K-l���A|]]�1�R�4�Qf�`�����^�k�R;'�b�/Qg��B��P�y9}Ռ�U�8|��ƒ��!O���XN�mo:Z }ܶ�'��Xùhe=�]9���v��!��G�*Q~�/?1{��d5��^ߊ~-q.T��� ��v��^I%By�؉h��Ew���C���^��`�[��.;��
���Η"��2G�#�3w�����uK�� s6۱w�u��t{v߽�_Xɜw�����۫2�����tP"<]��/V7�� �����n`n)>�0Ƨ\�Zoq���G6{6P�Uc��0�H\u٩�+���6�p4BḠ���q����PG�����o}3���*#Hsߣ��ӖG�s~�E3^=q~�k�Kz�����0�ҘC[��ra��� rs^��-�H�o,c]�U�����Ƙn`�| Q 51�[��{H����Ko����
w���Z�+#[RX�C����1��uJ�;���Su����c;�^ 3�������8;�?\�{��\���δ�����Jf���eu���n�.QuG��D޶��˖��3®���a�{��ԾtL��J����
���z�_¯R���ӽqb����m��@�'�[��� j�_uE����-��B���l��;�5a1�$p���`ݻ��ȧ�dX
�4&g���_k������ظ3�z�d��w���j'd�"S8��a�f����Va��c֍R��������L�&��?�^�A��Q����u�}�p��-|�8fJ��?�<�̛�))"� ���P����v(í�zF1��v����h�w��j�{F�>�H<{odX0�*�����L�~zb�04�R��B�xs���2+~�C��ٸ�ٸڇF��\��'8�E�o���Gw���ץ#�L�bv���<���/�u&�\���B//��{#��Wk��N��U�H��Mb��ɨA����G~�/�4�!�U�W��3��Rz��̺訩3\;�t.����r�ry�t�N��!2WC��]�l�Z��a�n�jј�S n��Q��ݺ��~V�Uhs�Ĕ��F�I3v��X�~�nVu�(�_ F셄�I�������B�j�k��wgM�����:>o��W����'DdU��M�����S1jw�3�9-1;-�Mf{��8�v�cԪ�M�^�_��\Dg��D�a�!��+Dz! �c�L�Ѧ��Gmv�ᇠ�|��>+x�U	�?z���S�//ص\�׫��FIfS{=E�_�n���Xb�GG�N4�rka��uU>iE/[���A��9�z=!|d�8F�xd�n��9�9l���ۧ��]b/VPs�iӈ-!�ᱵ��kH���a�Β��.x�����
�N�x28j�VF�ב.ro�@7��������S�ը9�4F�?I<�zm�=�"ボ�g�H�5hN�d���m%�ݫ�p�	o<��sn���D1|O)�<��e.�K�$��o��/��C%��!M�	,��1����-��Y˹>�V����Ok�NO�E�4�䲂���(>�I,��ʧ$����E�_o~}��d_HT-��l$y�,:�;C#s��ҳM="�-1Fι'�ᷬ7�LW�!O����~���gƩ���l<39!��	�ڗ�Z�)�j_X���0&��z�,7��-i|>�ܓ`�ZL�ո�!�����5j��:+ZΘJYp]V��o�Jyx��1'�.f/�]�?|��Sy=r�K��-l����xZ䖭�v�^d�+(]]/m��tQW?P��;
��K�|��r��"=��GIp����q�W�'O]8.kX�.&���ewt�6�*$0Ю�w# � -���̾�� �k������<�� )�W�a��3�~:�3����-*ymo��:g0jz��k�4Z�g-�.Gzn[mU-i.k��Y�]n���W6Y����
	���O4~'RN�LW�� ���\�ǧ��"j��d(c��9*���PM:e��瀎y�߂C�U?�OSݳ9hA.�4��!_�1p��g�-"�܄baw���}-:s��i�Ml��E���Pʰ���~���qn�	�)���&����+y%F��ᄸW�'5bP�M�T��uyB\�����]����V��#4��9�YM�uhq�9�#8.��cȂ���&�g0?�_�*(�+[{{D�o�>�4I�\u#ĭ���SY��Gۙ��k�g�`���{P{?4�_�kq�bg~㋱���g�6���%��~ւtE���Ok��q/��9Tf�JBq�t�����τ�ѳ�,6����WjQ��.Z~�0R��r=��(F	����H�(c
��k4�幨K֣F��i��Tz S�4�__'��̂�������r�΂���(P\)��7�I23WpZ̾�_̤\�Yy�3�Δ�t���ف�+�.��w�b�H���t�q��7f�
�|��:5Q�%�y�z^<��`vd�%��� ���Jf��h�w��H_���>͓i�� ��e���8$�J?�f���H����R]ge�J�v�D��r�ύ`2��=Y���'\1���1 ,J��d�e�(VDTK���7�#��N�������)�[R/�nNh�sz�&k���w��j������A����>7<������a����*���\ˍ��o00&�)���_<u`��	�B��GO�pvOP/���JLgA!�p65����q��������%o+�>�{j�������PK   ���X��D>  ?>  /   images/681693c6-5654-47c4-ac94-4786caa34b62.png?>���PNG

   IHDR   d   �   (�-F   	pHYs  ��  �����   tEXtSoftware www.inkscape.org��<  =�IDATx��}x�u�?3��ŢW�;ER%QT�:-Q�r��{�{lŶ�����;Q���ʲ;J,ٲ��%J�D�)���lߙy�3�X� � Rrx���3;3���Ϲ�����6Y�H���K��W�৯� �� M�m[�/���%���q�?�o\W�eeAܳw �n��-�Ć�����߄������x�=�]�q�N�<,|�
�ǎ^ܱ��H���P���ڃ�T��>�����R���`wW#㺤.���_�i�}^U���룿oD����?Z�C}1lk���4>�6���˱q� ��B'.^P�Ｅ^��?f�}�(j�eM9n{�	[[G��˪q��R�b{݁SʲqaM>��H��6 a����m�l.JJ'W/*�W���gj�ֶ(���Q�0zQ��T:GS��LbOw����͈���{����rܷߺ�߹��!�:2��܃=�yZ���,Ë�a������\���X+�m
��7�"����>�'���a���c�o�`4��ҧ&��2�no.�y]5�ws=��a���](Т��>��>75���o���\��է���������a��"L��B �[F��&�z��De�$�f`���\|��E��CMH�l��YA�r}:��Z|���jB�俄+CB�y!tE�1�?߱BQ�uK
q��-YC�5�i�]�.�h�U�|����P+H�_����&�;�� ?A���J�z�
|��fv��t6�ޟ�ׄ�$?�����������|��||c�Ɵ�=�5����|h4qW�*���6�qmF	���G���/ .綍��W��	!��en��6�]y;p]�>���<]����S��ѵ�������DU� ����s02�C��g-|���p˹e�������g!l~a�p����$��;+;q�M�CqYZ������Q��ޥ�]}
��l�[VUa�5�nx��!�m�{��p������0ޟ�7\}��}£�����ۼ�/����й�7�&\}ӧQ>o!ښw!��_H���~]8���y	oY^����,�� v�|?��6�߬w�+O���T�bx�9�t�z�u���EFP��O0��
�_������`+�]����	̫Y�ζ(|�5�Gె�����꺕���� ���W���/nT���#��G|f۲B��@"y�u�W_�Ҋ:un��uX��,�ۊ&}|B��ZKs��z��#�d[��f�ڷ�!te"�5�i�XTQ�kެ�)(����Ê֍��_M�[��ҳ.BE�bu��Ek�x�
,}��Z��F1,�uK?��P���7aϞ���GԨ i��{��4+/� �c ����ވ�ͿV N	2`�X�&,Yv��P�"З,=˷6a��P��h k.܀��buݚ��������t��f1��Den4<4�|<��e�sK�MJ8"ajB}�n��&Yjʄ}�lg�	yV<C2W��	ʳ|���,[�/�t�5���J]�-}
p�Ȩ�?v��K�L��H��5!�%!b*� �[0֧���aZT�p��g�}�w�)���F2���&�	d�4&���G۴ �Z�q��'��W����hܻ;ۇ��Z(Tm�T,��Q/'�b�3w��7��Ϗ][6b[�Vc!*B:bb}JV�~���pɵ�����a�y���a�XoGGLl�Va��G�W�QQj�����҅��:4y>��H��X��=�̔pf>vo} ���q�,KK�t�#�Jl
���;�K�Gx�OD����y����i�}�ī�Y��� 
6�Vqdk�v�j<��[�%8��/z%�����)�K^��8�AA��2�%��,y`$ea$n���[/%�+q��Pd<�6�%7`��ÿ�X���d�ȽG���|$;Dw�w7(E����(��"�����&���k�Ϣעg�,<p"����ǖ��V�����}Q���`�Ǹ�^A��:�B<��]f�ym5޲���	���[î~�fbj>�_�,'�N��н��El=����w"f��OEW���y�R����M�g�Z4���[^B����Rע9Y��^=�?�_x����FF���o'W�$/��ɸ~��C��,��|�)|�YQ�w�c���w_�I�u¼)D� �b��-�1,H��#-b�/��n�}m�I�\e��
����S1-��b���w�+���؛�J~GL�[]�O]T����_��_�\�7E,�K�"GP����u���	�*���u���O����5x�X��P�Y'\��w,�Ϸ�� G�/�Y���_F�F��Tb*,}�uy�xy5n���]<���*|��P�f1Ɠ"�Đ���ը-��C�k��lӻq��A�JhWq�޾���bp������B1�I��s?|�B\/�m8�(+[�U���v1��"f1mn��o�P�va�4��u�ů 2����J) ��-E�x|uѢ����}Gā��֍G��7/ă�D���|4������GZ���m��lX��pRܱ�/�'���R������o߿D8t�O��hRN�m=��1d�C��>�����m6cT�r�b��Ou�5�h�i
��kg/~(�mȟ=2�F��P�`,%�u�~w���qyM9M���A��K���k�*/�Q�~�S�hPy��x]����hJ]IXʳ'G�	�}
!�A���^�����I��}���#quۏ�u���!E�v�u��I�>�%p3�����q�Kyݾ�(>p�a�����$�bB ��t�1-���e�Fz��!�y���`�PSf��߼�|C-���^�����Lѧ6�gO$��p��g��rC� ��>Ǯ#a��)���<���I8�"=��S�C++��.۟��Ag1�l�<|��u�'a1C�Oڦ��3mn����Z!TJI�	�Ol41����&k�i�7�"�27�sK�	�ØM��o&����/�;��9n
!I[Ǌ�!|��&�-��@���0O2C��M����芕�P��h6�q��;ѧ>����o
ꎃG�9���>�rs���4)�N� 	�\��W'ě�g�6�R�ki���k��I<�>��ӌ��ަ�(N�l��(,Y
� ���JA�S��?��]�M	��u`�у�f9V}�nV�b�(�K�c���O-��<�Z����Tr1��7���u��4�P?�s�1fF�4��V�P]~nB99j�9�"�D\�4�g�jB���p�h�|�BL_/�z?L1<�i�>�!31� �TH}ک^��Q����S>h2';'�?��L���RB�<3�^|6M!��-�G�w��<�'0�8Y]�|�DW�1Rם�&V����|�Zl�1�r�E�"�r��O�Y?��/�)��O>s�
rst�KnAϊ����969c^��]��(ׇ��a��\}�C��
!\n����H�}�twU.�&�\�^C;�<"@��F��"����tw�'sޱ�#N��g.9�f��@�f�����!������̜T݇���c"K��D�1n��y�5�$��i�N�Q;��=�S��^I�R(��Wˮ�4��J��u�=Iy�֗��M87E���644�Dr)#'cٵq�:��4�"���7d���K�:��2�! 9I�h�̈́�x�_���>+��r�ײD,������Y&S>W�O�Vݸ¿���*������9�"�%�){*���x�g@��Y��/��c��wc�]���H&x�;ߊ��K���� �^W��'k{q�]w�A��/++ŵ��>�9���5c'��p�9/R@%�n�0������s�0����AH�7.���?�H$� LĿ�������@_��=����J�Al��B���X]Bii	��[P�O O�*WK�di!P9��Dm���E\͛��d?a; ��,6�#�IB!8i�K��;��'Ї�s�g6<����E��]
��s�X*��v�8���\|��O�8h`0Ǔ[��x�I�\�
����^���$�`$U��@}�J���̿��yf��L��4���k����-7Ll|������h�r]<1RRf*�%C�`�I,��c��DLh��-�����iCi�����[<�қ1�v}����n��⊍ruOo_�o��$#z�D��'%��]V� b��!>)*�� Em� ���Y���1T�ּ1}�eSLL��1�}��]�cV�fFyY��5*V�Z��#��(��8,��!�J;P��t�ir�7�?	��.��".bӢ�5>)(�[�<7�坐C<��	A/X>��"�|�䖧2f�Ī�Y������2���C���˗�I5�e�I�,���>��#ibT�S6f�\�S��0��(�8��z��N��23m����K�8S�*�R�H�$(��d�>$������"�D��V�Àf�H����s�z�ODD�^�-P�)'l�G���R`pUy)"9�hL�)�ז5�ׇq�����P0�E�cǠ������&�p�,�nj*�8{b���ߜ�^�#� ���ڢj�n���◝�t	�Gr0��f)c~�@���}~3^���8f�����T\�zi�>�{�,+Kt�I�Q�������\�b�����񛿄����x0�=X�>�*�G�>�E!���Q��ڑ4�D))$�� ��ea|��w"�`������Ư��ʰo�L|O�?�����9C��@;�'����.�}Ǆ���b~]bb�����N&�J��ʠ[��!~���A�rJV��1���B�WU�$FOw�*�p�D��.'�ru�v~���G�1|��a�~d+�Ǭ,z�@��á*�~�|I����q�?�6���gPG�U�����)*).�֣�%3$�L�_���2�T�oSot!��B3�O�������Z�"ĺ�
9��
�D��c�L?%C���P��ʪą@��Y�ɢ�BS�_��d��sޜ���A�pL��1G��r����Ю��;�E(h�az�3�l�)�����$g ��j�V:Ru�<!2�/{c6�z��%���?��0D�O�~����$���4r�B�AX�Ō���+͘p��N�����a�ј9M�n1%�Z��a�f����b�-�5`�Y�v� ;�5a�l�oj {�?�H���9^������sވx���8v|P����Б�*��/~�Z��!;2]�P�$�I�� J������?��ؙ�"�!�8��ԩ�h��˜����b�מ2�=��Ԧ����̞d���B9/��D8��?֯_�b�!ñ6��5����� FlACc���L�k�C{�Y��p4h^��̇���'�N�,����.cbIk�U*�G�`^n���m&�A���ƺ^9�'�<[S�V��D6��>P3�{�W-���@ ��������B��v���9�^z�c�D
�ΰ�qg�o�ch�� ����	(?dCQ=���xC�B̻��S��yQ��2-��jq}�����"8��RN,'9��{tM���oR'�Q�P��a4Z%X.��^����kUb�ރb�3ڕa����#�eH�8'��9�B6Mž:�W��+zȱ:�C�DpU�[�@�����VN��m|m�h:�'�Чh���d�=��c�4��v��$�M9�h�Zu���\�Ԉ��/��M�b��S�Q��pj�5�R�Q/T�/��ADcLr� �T�6L��'SɄ_y���3��t�$�]i�PGܳoV��u7�W�s�38��rǮ�������}�oN��C�·6w��Zx���l���zm�pF���D���>q�"f=��\<l.��<�I��s�|�p��X�<��ʩ���4���F$D�)+����,�O����1�Hg� �χ=�Pk��Β	z-���M��訍_�T���:�e?�]I���x#@�S����6��g�JS���N��G���H�8Q�=a�n�������"�����m:���t˩5�(i�`��b�%!�X���Z`~�K=�ŵ���k��R�5�b�7����F {~É>}�gڔg�=#�K��&�I�H����BW���ocK��2a2%�8�0TpAA߸��ԕ+��VC� ��y����tI��n��m�c��z��n��*�H庖�Ѣ�]A�_�|��+?����=��+)�,#��ǅ�ˌ8�����cݝ_6�)l�Ϳ9����n������:���@�>)�s�8��`4�k� ����'B
w���R_�aw����2|z^����ӥ�i�p_�kꃂ�E��K�j�Εa��� ,��U����w��]��PQQ�?�)|�8�������Q����-�s����yJ���m�����&��\K$�tA�%�㐑n� >r�"�d�&50�YV]GU-�.�NUO,�,�5P�V,LS�X�GI.�B#$JC>Ya��ExA=����˔:�A?�+K����8��b5�ŕ���>~�1�.fm�p4�$��&��b�gOmc$iT��MmL=�/:�}�#2��	�'BGR��WL~�`�D�<V�|;<$@�ca�9GC1��;��:���z��dO"+>����=τ��^�F�Z����>��;�o�o�0�O��������v�����&��w�����D�ﮰ�SÝ�\����Z_$�O�߄��Ѵ����΃�zƠ�ht8z�-��;�9�vv������X\��/��	��϶��av|���l�q���;�Z��pT�S3H��Q��4Co�v�s�4��}����Ǖ��/����a�M�'�$�)=�$~(X%��hW{�a�)od ���\����ҏp��c�n:!^��Z��s*u�hg�0���-�&b���qaNu��9�\��
�{���Ԇ�i3k�ge���j<�,z
�?�RW��y�*Kh��j��A�����8�-�o*y�,�����\R��s�)d���ˢ
��֧~|C�
��3��XW$�����Y	���7���}��(
jxZ8�p�`��Ѥ�m��V���Z������+D���b��AΞK}���ۈ$m������f�����5����)�����j/
īX-�a4aco���i�Q�4��*�q��H��"b�K>��L��yȑAK))C�b��2�~�s������d ~�=tRq�{4��S�M41�n2O%��{�L��&�s�EE:�_�����E��g	#���L�	�.$qϵaC�!pk��6����zC=|(ncG��t���R��s��X���y�e�AQrHwvD�v�X�q���ɅE�mn���s����AT��{��ykX;�=�gy���s��cخ
j4T�bs���H/�O�]�(��2]Z��&��Ԍ��-:���	Ǻ"R�%D�&�!�/�)�gT ��!����&��z�==��=`_�D�ʪr�YGGt��q8	81�����7�wb}e�e�Z�h�B��	|���?��%U��/Oq��rϕI���-)4�^-DMvOJ�ab��a|�r���C��j-Q���E�g�m*����/��a�r����]A}��HSz��A���(\A��ȡ�!�A���}x�1��;��P""O��C��8�T��.�=�!���,�(s8e�tB��O0�rv��L��?���m���u7�W�De�t����~+��� ���:�Ƣy�1�i��=���z��8U�v�ݏ�<��o[�J���P���w⎧~���G�kQt�`yr�����PW�T'��Y`D�3�2A�N�Q<]\#��d��VS��Ǵb���m�	�u��y��*!��4���U�w��8r�D������h��9 s�l/|G�O��ǯ	�>�K��2�x�m�{2�E�I��w��&XPU��V�1'j^���M�5u�C�t�vFhJ���7��v�O�V=�B��WҎ	PfWH=Uʋ�pѰ��
Ȫ�E��!�4�ISe:��@�ꛓi:���8��@ �J_�	�����g3�v��椒2�<��we�݉c���ZR��[e��jqi
�@wa��h
�)��$w�j���Y�s�C@o�J��J��r�;�˰4�:s�rm�ǚ���4l��N����UY^.�k�����\g��)�U_A~��,Q\���҈��	`ѢE�$�R���=�d���k�z��\�%�O`�h��Ԝm;<��mV7��� ��v�U���ը^yeV[Jq]qI).���*,�1��9&T���q�57�yN��mC0;R����I��g��R���q��KǛF`��QYQ]�7��3J����"Y�����#l�<Vxм���Nۮ�d��w$���BZ�/]D�?I_����z�櫉�N���'��}X��G[=17�I�kb���Q�%�4c�]�m���e���H����h���6�=����f�r�U�or�{�e�!1��Cfڴc�L�[��Ox�v��NQ��SiDؙǎQsf#�S��:c:x����{�������:ӎߴ����9Ӳo�:$�!�BNe��DV:�z�C�����0�������v<�׳�� �7o��t��K3� �4�t+C�x�"��Xy#5o�|6��,�{��O�R��Jr4�.�Fj�AM-����A
�ׁ�K*cJ�znL!������m���v��F-�<{�aym<�80�N���eN�=�[���"�By��z=��ziF\�~��ě�j�/3j&�YNM�xJ�O�RW���:��L����U�kX/�G�^WU���r�d"�y�Id����c�Z;���2�
?�}p��9HL�p�'���:��Wj�^��\7��d2 �5����
a�SEH�%BXL��k�f"��D��T�DdqAhe��2+�I�Mgc�y�R΂?�yU��i��^�3D�v8	m���b�H$	�CnZ�S����'�%* ڸ���!��T,*�r�T�~�F!��)Lv9�t��\Q<�LW��ϴ���^<j�A ESxhR�\0��e����1S��~����9A��V.���uRr��iX)�&u1�Z#��)�p�ٹƴ�NE�24�u��
'͓ ��+��3�:l���C�O��y�7ݖ�D=qs&�8AV]Ѳ"Փh��/�F��I�-(d*��-m&��8��:��I����<��"���d��\q�g��,���<�$saKqs�Y�A�BΟ.�d&���{�d?&�J!k��,zL�1�\�a2�i�J#h����N�ua�m��=�Q�ٽ��r�7�Rp��A��>M���Q[���ݖ���_f*�t�S1-{�L�!i+��}V���
�i��1WO�Xw��&3I�\���1����.�ud3�uo���/�m����P4DW����XK��4ԫ��#�c�<�)N1�R�.����O��%<O�we��Rf9'"���0`)r:\�L�L2A���U7К��eG��
�暽�r᠝2qN���ɱ�������EL���x@5-[�ɯ,b����|r��7y���t�a ��}1������9f�3�s� �O���1i��Ǐ�\g�RB�E""��L.f�,Eke���=�#d2�Ho�鞛]�%_ �AJ�gˁR��"�R��ĸT�+�h�Pw<�2fyёd�Q�3���9�x~*�|
q���!S�n��CrsI���|?j��s��-,}��H#�Ф����� �>5���Q�B������wY�D�E��1j��wf�OD�bXs�*q僢6:R��E�W��4ʤ����g�L)>�V��ZG�QD��
�"A+����U[R�Mބ89����VV�q�B�v��J�SD߇���ŮO��6
�P�6;ʛ\q�<��t	q� � ǩ k��^Z����Ŗ6Ag&[{m�b�^8)���b��$b��sj)<qV)ȣb}�)��g��ٮ�B3�I��q� 㒺|����Q��:���2��L�,ۇꯡ$���c]MH]�rۨ�~0�J0S�J�����E�>�����1��j("�;b	W��s�{8+4���2EU���U���"@�}8���G�cǬu�*�E�-����e�N���>����/���<��g���PL鄩^�̳�o�dTXb��"\P��A�+��5˅�m�{ЍSqL4.X����� �PLq�Dȁ~��(�V.D�8����4�dr�\9��k6E:��I��$����3:Y:�ku�1G�QܱP�ѕѼ߯�JL�=X<d�;�1oymO$�g�Fpò"��g��$�6R�cx2z��M�)��@�&�Ϸ?@�k+D���5J�X� ,��Enp�	���B��R4E���Gt����58��XC��:Ǵ�X'���%y�8���ܱ�<U��Z��#:�}����犕��쿂1v��Ek�i�$n�D�D�p޿�&g�n���~��Jr��^���:z%A]�G�� � V(���K[H|Ur/7�<ѫ
'[��R�^0+�8p��#I�5/J"[�D^��p�]1$e�3F\����(8I�?�\�TL["��Έ�X������e�6�]�OR2p���P�:{[��}=1�U�g�`wWT=/��*"l�CQ�#q4Ct�Kh<��h�Šj	Y�ϗL���3��tp1�Ef�Cl��ܫ;䱪���ci,z���q��<YߡJ�/�m���|"Ǔb�%UM][��Ӎ#h�J�Y�)�V��:�7-�QKq�J���yb�qs�R��M���GY�ٔ��c�1Mn�G�K��s�:A�˩Nv�ɹp��i'�-�g�K1n�5�t8�w<� U��[��c8�W@J��Mм�v�SH���j�yi���\�E%9��$���Y)�O����)�2JP��y�_WN)�+.jq��Q+�a���HH<Jlڎ� ��ߦ�ټz��"f"-sm}֭,O�yΜ'F�u�rNF�Gs�Sn�#c}��ջv�N��bAE�"�"�V��wμ\<rh�Ą70�N�4u��+aE��%��<���ǡ�r�t�`�c�q�Ǘ�f��w���1|'���D�S�b�]id6��F�t"n(�#C)��y��� @����pS��G06���Ή���r�RǱ+���*�Is�C�T�O�ҁC�5|良���F�QSq�����Ն�^���S4�t4��*�	���s����Y�D���W-�w-&o���-6ƊZMkl�����|��hV�~<�C�M�M����M�N��U�&��QtȜ'Z<4�� Ԩgt��ꍕ"��^T��Z:y�-�6�q� �k�S�Җ��/�?+�v�����c�+��p��
X�9�#ӛ�$�g���Z��>v��p��L�s�T�(���o;'*H��4�nB_$���vx̤��(3��C�|M<�8���]+K�v�]by	lDFe�S�~�x弿Wt����;�MX�d�KZw|��e�'�C�&$0��<�7D𞨋 �E�(df��v�5.Ff]d9�P���1������Ds���C��&r)����V8 r6���WWW�b��Q��("��N|���V��B�3�!aE���	���(���(?�A�p�T�X����A @�p��*V�9�D9�9v����0.��shg=�΁r�� ��"�����NiN�3P<2�8��F��GM�!#r��I稩�2w���[oI "��=s��t��c���\���}'R�3�$Rw�����m�=�L�{#�#gcl��ɋ�1ǌ�K�\�&�$��r�5�?{¹9Q�CU�ND�"����8�$��㤽X���}W�s�5Ǝ����8�t��\%��;oS�P��ꓙ&��t�Cd�W�CI3�������&',+uV)��ȭܧ�;�,�$�ވ���c������6#�3M"�'|�ͪBQD�S,1Q�S&wV�Oq�Di/+�9bI��Z^�Sg� �g�jWT�F��)�B�K�T��y�������CD�sD����S!:���/�]����䲑2y��L'j0��r���L��sH��5a=���F��R�e���
*>�q!RS��/#���\�8A���f� �d.1y���u
��{Z��@�&Q
����?���1���*��v6|�)�c��9&9."���=�\��B�k]N���:?C��U_� �+�l���I��r�B���6��f��=��1��+��@�CS�������K\�Y]�E('�ͭS�[�S��Nl�8�H��!��g)T��4��A6�r^�M��8�U>g�a��T�;�˼�C4LΣ���.�r��Tnju�u^Vb��4ƨV��.�A���d�$8�x:-ST͹�N����bל$����b����F7�cE��|�Ikݼ�����&��B�l��+�^��L���$ }�T�л��^���:���"�吺ʔ���R������F�)�8c:,�צ3��I.��M"Ӧ�>':���&��?8�^���cҮ�Xu(�ܱ��@����M��Kk<��&�����2g��U���c8�\A_�B�gd7�r�/�|U�J`�j��r�CYk�:SN@��e���#��*���?a�uF�p>�r��Nv�N�2B<�Ek�J��f{��}*�J.!�Ѽe:�ܦ��2������S%�9�'�E/|Py�cps�|S@�g��	gb�WnL�e�0I��Q��4�i}����;t`��ϝF��Dz'�s*�8Y�WS,Ѭ���p�J�kEC�q3anɤ^CNbZN8�}����309����>�:��aV̳-f�f�	uE���I��.��gPQ5Itq�YGIg��M\�$��A$ЙM�M�_uu?/�6x]�+"f �5ӵ���Q�p�W���!�7��ʞDD�q�%	��8�p����� f�1%�2�43�D@.Qi�}Nu��NG9��Fky&�wv;��J�ce�i��ƴ��P~C-3�d��Y�}b'����l�>17�M�>��P-*/�}���Y��X*	U�C�a�+�G�cU���4���ݦ0��!lTv���(���'�K*���=��R>��X6���袧�T[*��Y���)3A�X��)\1d?,�a��^��,�w���0��^'���E{�#n�ZAE+�����>�vJ8�����z�7WP&S�Ӿ��R<��R_��Ϥk��<��&�TYt�Y��e���z�}�F���ey���	���5ϫ�`}��7=dL��P֩�t'2�P���0}��44ϫ��01c�1񙓝;mY'T�odx͋<�֐���)E�	^��!�v�~�e4�xf����i'nSI���!L�qvR���ʛټ��:�d�g6�}&����x/�"�N2����X��
u�N3�b�ݎ��fI�;nF��+����Dj�Y�S�c+}(W��c�Z�����,�3�����}�U���ѱ5Ь�e�����5�ډ�2KR
����I��5�:�(���LΒ��o�p0�`��NOXR�B�'�SX�o�4��Q��O��y�:�vS�B 3����ދ?�x޵�De�on�Ç�������O��޹X�>�\G���mNb�'�"�/+�W�עs$�����ZT)�?o��Ҳ�Ԏ�~��w�g�Bl�x��y�o^\��\2O!���_��>��o_Y�����ُ;^�QH���$�s�>�G�I��8�R�~�6B�^���ksp��R�r�%TV�7v�Л��w��%�[76�,�x�|�jg
�;n�܉��է�qY�Ƥ6����m�~��* ���*͔!g1�+O��޳T��
��C�L�#gy�/���ۨ�~�X.|�a�)��������}N�$s����� Mu�y'�h�y�K�:��7.��I12�0�\���o�Kp��K���o�FQVЄ[����_��ԃ821W�f�%��"4�Ǖ(��<�L��܅���Fݟ���n��m����D���W�êP���?~�"l�?��)J�)�8^O1ű'��B��_j힥����e(�ĥ�������W����w��l�,��w/���.�'M�՟��^��:���&���&6���P�߾P%��գ�0M'�����
��=�*�g"H��xa25S|X�I@���RE��3G���U9���mQ|Pg}�6����G��j]���S"2���"�&��Ay��/���:9��Ib&�Q���j22�g�7E�p̔Ɓ;�+uK���E�E��t?։{��s��~r\���M�6��x�[��M6��>�)���1��<�>Ӏn ޻o@�R��EG|�:T�����l[%Y?xpI��E?�j��������{Dq
E$�p�菜I�����JI����|*U�D�l"7�B,�o�������v��J�_�����_�E"�9A*рOOo���VP(��T�g����bi����)*�+b�Q��XS�RN?x^9^hUȾ�*{Y��cD7�N���~,���xE5��X���#��gu)>q_�B�gO����`O���l��c%	cgg����-dr�����d�"�ơ㚊�"�8R�CB���I�)��N����$���[*q��P���*��xn8n�<,CD���W��[�T	�o߿L=����̯����O=� �C��j��G���fU�N��ߥO*�|�Emh3Q9���g���˰�����7ԙ5��
���dm�/k��]W��U9�9_�����F�F�����c׿{�MM���\��nb�g^2��_D!�}��Fu�5,#�=�0g��±�:�~�_	 Y���OE]��ͬS'`���#J�(ȉ�W��LGr�i�K���i�q9	ݓ)c��o��5�
���lD֗oU�3ǭ!a�0ӎ���"ޓ<wR�x�2{�a�����٦���?<ێ��ܲ��W�s{�hVb�xm���i��3�9oOs�#uzf�T��[�55�K۸�6�w�"��$m��xjl2]sj\��M֜=SRx�V����Y4�wwG������h�09&r�L��3��YZY^9W���NS�M2Փ����~�w ��7�(<�&�Қ�\�����@��>�s�)K��[�����3ճ&S��-�p�3J��B�D�h�T�P�y�D�ԍ�v�J$�|a^1���W�+�T�����Ɯ)n�}������39#cR��BF>O���@1!-���֜����[3aA�e�)��_81��Q�b� 3z�hl>�i}p���v:B2ݓY�\�$���`��?��+sN*.a�6��^��8A���`v$�Z.�ᆚNQ,� Yv�=!��gU�T���d0&@3��Y����u���@�b���EB��Y������k6kcXf�d�;,%�X��0`N�C&�q77�2c�Il����l{�)VÊ2Mm��}9xn��F�6�-F��,�c�1�2��B��$h�{�Ddn*L�9U��L��@˄+����\��ؘ��N���f�EW��8N��`:-+"����SK��}Y���49x*y��!p	�P+�R�������csӎ���-�BB92�Y��Nuc����2�c��0�6�����lSz�[�MA�yZ(�cL�Ζ��z�Ck��&�0M�������i�\��������2��\    IEND�B`�PK   �N�X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   �N�XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   O�X��?��  5     jsons/user_defined.json���n�8�_�еi�(R��val��Mn���(* K�� �^Jr��]�w2E~C�����Z��ou�-�Y^�4X�u��Ui^�%\"3���0�V_�_\�ð6n�>/��W[3Q�N�U͓�\檩TUvMU�	nc��1�*�E�AnL҄QH gN������8��mkݪ&��i�o������(Nd) �G��(��p�C�(fJ�e]ޙu�C2��+��Y�ee^�y�)�*X=eX�m]ȧ��h��FKf�����qM�S����7;*7�kr��0�j�a�yaFap���"o�R�W�Y���7GS�D��������b�l,��������>~rb��e^؝nu��zaɒ�8�Ԧr/*s3��^̿��VhC���C/�sA��^�:���t(�w&r��-+��1vCmQa�쏉jK
��~L�P[P�/�c��z�"�������g7uFQ�����M!?l|� "[V�qO���B��F'�����X��̥�|�n��K+�ź�����'6rSg�,�In����j�P��jk#Oj��/�����{�xR��\\ԓ�����'խ.2sw��T������=�F[�c�e��yc���ʴ�S��BRA0P�Q@��@BDbz�$������`�MU�ˏ���7�i����<ġ.�!�~tf�0�|[wl���myQ�;��M��I��5���;6���"ʲϤ����_BOF�m�P�%U�����O!s�y�?W�'M�0��7%ս����j�i��6��_�զ���rT�k�P!1�% b��@�4I�R*�J�*E��� 4�
$� SՄ��g���%I(L='*,��+
���'*)	MB���ę��b.	�cR[v�%�Si�Kn>-L�4���A;ٝX|>�1D����>ç�S ��\n��3,�"p|F��~{�}�S�(���{��#c �C� ��:<`�?�n����� ��<�|�W�g�~�}�PK
   O�XH���
  AW                   cirkitFile.jsonPK
   ���X� ��! �3 /             �
  images/199a26a2-2ca8-4fec-b52d-fcf4e34cacf1.pngPK
   ���X��D>  ?>  /             �, images/681693c6-5654-47c4-ac94-4786caa34b62.pngPK
   �N�X$7h�!  �!  /             �k images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   �N�XP��/�  ǽ  /             Ѝ images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   O�X��?��  5               "@ jsons/user_defined.jsonPK      �  QD   